module rvclkhdr(
  output  io_l1clk,
  input   io_clk,
  input   io_en,
  input   io_scan_mode
);
  wire  clkhdr_Q; // @[el2_lib.scala 474:26]
  wire  clkhdr_CK; // @[el2_lib.scala 474:26]
  wire  clkhdr_EN; // @[el2_lib.scala 474:26]
  wire  clkhdr_SE; // @[el2_lib.scala 474:26]
  gated_latch clkhdr ( // @[el2_lib.scala 474:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign io_l1clk = clkhdr_Q; // @[el2_lib.scala 475:14]
  assign clkhdr_CK = io_clk; // @[el2_lib.scala 476:18]
  assign clkhdr_EN = io_en; // @[el2_lib.scala 477:18]
  assign clkhdr_SE = io_scan_mode; // @[el2_lib.scala 478:18]
endmodule
module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [95:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [63:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [63:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_scan_mode; // @[el2_lib.scala 483:22]
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 187:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 323:36]
  wire  _T_319 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 324:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_319; // @[el2_ifu_mem_ctl.scala 324:42]
  wire  _T = io_ifc_fetch_req_bf_raw | ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 188:53]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 255:30]
  wire  _T_1 = _T | miss_pending; // @[el2_ifu_mem_ctl.scala 188:71]
  wire  _T_2 = _T_1 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 188:86]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 553:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_319; // @[el2_ifu_mem_ctl.scala 555:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 189:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 310:63]
  wire [4:0] _GEN_437 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 671:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_437 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 671:53]
  wire [1:0] _GEN_438 = {{1'd0}, _T_319}; // @[el2_ifu_mem_ctl.scala 674:91]
  wire [1:0] _T_3079 = ic_fetch_val_shift_right[3:2] & _GEN_438; // @[el2_ifu_mem_ctl.scala 674:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 325:60]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 277:46]
  wire [1:0] _GEN_439 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 674:113]
  wire [1:0] _T_3080 = _T_3079 & _GEN_439; // @[el2_ifu_mem_ctl.scala 674:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 660:59]
  wire [1:0] _GEN_440 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 674:130]
  wire [1:0] _T_3081 = _T_3080 | _GEN_440; // @[el2_ifu_mem_ctl.scala 674:130]
  wire  _T_3082 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 674:154]
  wire [1:0] _GEN_441 = {{1'd0}, _T_3082}; // @[el2_ifu_mem_ctl.scala 674:152]
  wire [1:0] _T_3083 = _T_3081 & _GEN_441; // @[el2_ifu_mem_ctl.scala 674:152]
  wire [1:0] _T_3072 = ic_fetch_val_shift_right[1:0] & _GEN_438; // @[el2_ifu_mem_ctl.scala 674:91]
  wire [1:0] _T_3073 = _T_3072 & _GEN_439; // @[el2_ifu_mem_ctl.scala 674:113]
  wire [1:0] _T_3074 = _T_3073 | _GEN_440; // @[el2_ifu_mem_ctl.scala 674:130]
  wire [1:0] _T_3076 = _T_3074 & _GEN_441; // @[el2_ifu_mem_ctl.scala 674:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3083,_T_3076}; // @[Cat.scala 29:58]
  wire  _T_3183 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 333:30]
  wire  _T_3184 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 333:44]
  wire  _T_3185 = _T_3183 ^ _T_3184; // @[el2_lib.scala 333:35]
  wire [5:0] _T_3193 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 333:76]
  wire  _T_3194 = ^_T_3193; // @[el2_lib.scala 333:83]
  wire  _T_3195 = io_iccm_rd_data_ecc[37] ^ _T_3194; // @[el2_lib.scala 333:71]
  wire [6:0] _T_3202 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 333:103]
  wire [14:0] _T_3210 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3202}; // @[el2_lib.scala 333:103]
  wire  _T_3211 = ^_T_3210; // @[el2_lib.scala 333:110]
  wire  _T_3212 = io_iccm_rd_data_ecc[36] ^ _T_3211; // @[el2_lib.scala 333:98]
  wire [6:0] _T_3219 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 333:130]
  wire [14:0] _T_3227 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3219}; // @[el2_lib.scala 333:130]
  wire  _T_3228 = ^_T_3227; // @[el2_lib.scala 333:137]
  wire  _T_3229 = io_iccm_rd_data_ecc[35] ^ _T_3228; // @[el2_lib.scala 333:125]
  wire [8:0] _T_3238 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 333:157]
  wire [17:0] _T_3247 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3238}; // @[el2_lib.scala 333:157]
  wire  _T_3248 = ^_T_3247; // @[el2_lib.scala 333:164]
  wire  _T_3249 = io_iccm_rd_data_ecc[34] ^ _T_3248; // @[el2_lib.scala 333:152]
  wire [8:0] _T_3258 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 333:184]
  wire [17:0] _T_3267 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3258}; // @[el2_lib.scala 333:184]
  wire  _T_3268 = ^_T_3267; // @[el2_lib.scala 333:191]
  wire  _T_3269 = io_iccm_rd_data_ecc[33] ^ _T_3268; // @[el2_lib.scala 333:179]
  wire [8:0] _T_3278 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 333:211]
  wire [17:0] _T_3287 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3278}; // @[el2_lib.scala 333:211]
  wire  _T_3288 = ^_T_3287; // @[el2_lib.scala 333:218]
  wire  _T_3289 = io_iccm_rd_data_ecc[32] ^ _T_3288; // @[el2_lib.scala 333:206]
  wire [6:0] _T_3295 = {_T_3185,_T_3195,_T_3212,_T_3229,_T_3249,_T_3269,_T_3289}; // @[Cat.scala 29:58]
  wire  _T_3296 = _T_3295 != 7'h0; // @[el2_lib.scala 334:44]
  wire  _T_3297 = iccm_ecc_word_enable[0] & _T_3296; // @[el2_lib.scala 334:32]
  wire  _T_3299 = _T_3297 & _T_3295[6]; // @[el2_lib.scala 334:53]
  wire  _T_3568 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 333:30]
  wire  _T_3569 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 333:44]
  wire  _T_3570 = _T_3568 ^ _T_3569; // @[el2_lib.scala 333:35]
  wire [5:0] _T_3578 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 333:76]
  wire  _T_3579 = ^_T_3578; // @[el2_lib.scala 333:83]
  wire  _T_3580 = io_iccm_rd_data_ecc[76] ^ _T_3579; // @[el2_lib.scala 333:71]
  wire [6:0] _T_3587 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 333:103]
  wire [14:0] _T_3595 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3587}; // @[el2_lib.scala 333:103]
  wire  _T_3596 = ^_T_3595; // @[el2_lib.scala 333:110]
  wire  _T_3597 = io_iccm_rd_data_ecc[75] ^ _T_3596; // @[el2_lib.scala 333:98]
  wire [6:0] _T_3604 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 333:130]
  wire [14:0] _T_3612 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3604}; // @[el2_lib.scala 333:130]
  wire  _T_3613 = ^_T_3612; // @[el2_lib.scala 333:137]
  wire  _T_3614 = io_iccm_rd_data_ecc[74] ^ _T_3613; // @[el2_lib.scala 333:125]
  wire [8:0] _T_3623 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 333:157]
  wire [17:0] _T_3632 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3623}; // @[el2_lib.scala 333:157]
  wire  _T_3633 = ^_T_3632; // @[el2_lib.scala 333:164]
  wire  _T_3634 = io_iccm_rd_data_ecc[73] ^ _T_3633; // @[el2_lib.scala 333:152]
  wire [8:0] _T_3643 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 333:184]
  wire [17:0] _T_3652 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3643}; // @[el2_lib.scala 333:184]
  wire  _T_3653 = ^_T_3652; // @[el2_lib.scala 333:191]
  wire  _T_3654 = io_iccm_rd_data_ecc[72] ^ _T_3653; // @[el2_lib.scala 333:179]
  wire [8:0] _T_3663 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 333:211]
  wire [17:0] _T_3672 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3663}; // @[el2_lib.scala 333:211]
  wire  _T_3673 = ^_T_3672; // @[el2_lib.scala 333:218]
  wire  _T_3674 = io_iccm_rd_data_ecc[71] ^ _T_3673; // @[el2_lib.scala 333:206]
  wire [6:0] _T_3680 = {_T_3570,_T_3580,_T_3597,_T_3614,_T_3634,_T_3654,_T_3674}; // @[Cat.scala 29:58]
  wire  _T_3681 = _T_3680 != 7'h0; // @[el2_lib.scala 334:44]
  wire  _T_3682 = iccm_ecc_word_enable[1] & _T_3681; // @[el2_lib.scala 334:32]
  wire  _T_3684 = _T_3682 & _T_3680[6]; // @[el2_lib.scala 334:53]
  wire [1:0] iccm_single_ecc_error = {_T_3299,_T_3684}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 192:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 637:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 193:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 194:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 480:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 194:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 194:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 194:72]
  wire  _T_2476 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2481 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2501 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 530:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 393:42]
  wire  _T_2503 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 530:79]
  wire  _T_2504 = _T_2501 | _T_2503; // @[el2_ifu_mem_ctl.scala 530:56]
  wire  _T_2505 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 530:122]
  wire  _T_2506 = ~_T_2505; // @[el2_ifu_mem_ctl.scala 530:101]
  wire  _T_2507 = _T_2504 & _T_2506; // @[el2_ifu_mem_ctl.scala 530:99]
  wire  _T_2508 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2522 = io_ifu_fetch_val[0] & _T_319; // @[el2_ifu_mem_ctl.scala 537:45]
  wire  _T_2523 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 537:69]
  wire  _T_2524 = _T_2522 & _T_2523; // @[el2_ifu_mem_ctl.scala 537:67]
  wire  _T_2525 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_2508 ? _T_2524 : _T_2525; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2481 ? _T_2507 : _GEN_38; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2476 ? 1'h0 : _GEN_42; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 194:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 196:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 196:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 285:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 285:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 706:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 285:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 276:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 276:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 327:71]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 276:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 276:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 285:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 285:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 285:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 285:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 285:114]
  reg  ifu_bus_rvalid_unq_ff; // @[el2_ifu_mem_ctl.scala 580:56]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 552:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 594:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 621:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 312:62]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 602:56]
  wire  _T_2622 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 619:69]
  wire  _T_2623 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 619:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2622 : _T_2623; // @[el2_ifu_mem_ctl.scala 619:28]
  wire  _T_2574 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 598:68]
  wire  _T_2575 = ic_act_miss_f | _T_2574; // @[el2_ifu_mem_ctl.scala 598:48]
  wire  bus_reset_data_beat_cnt = _T_2575 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 598:91]
  wire  _T_2571 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 597:50]
  wire  _T_2572 = bus_ifu_wr_en_ff & _T_2571; // @[el2_ifu_mem_ctl.scala 597:48]
  wire  _T_2573 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 597:72]
  wire  bus_inc_data_beat_cnt = _T_2572 & _T_2573; // @[el2_ifu_mem_ctl.scala 597:70]
  wire [2:0] _T_2579 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 601:115]
  wire [2:0] _T_2581 = bus_inc_data_beat_cnt ? _T_2579 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2576 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 599:32]
  wire  _T_2577 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 599:57]
  wire  bus_hold_data_beat_cnt = _T_2576 & _T_2577; // @[el2_ifu_mem_ctl.scala 599:55]
  wire [2:0] _T_2582 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2581 | _T_2582; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 196:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 196:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 197:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 196:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 197:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_319; // @[el2_ifu_mem_ctl.scala 203:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 203:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 430:45]
  wire  _T_2106 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 451:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 407:60]
  wire  _T_2137 = _T_2106 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2110 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2138 = _T_2110 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2145 = _T_2137 | _T_2138; // @[Mux.scala 27:72]
  wire  _T_2114 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2139 = _T_2114 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2146 = _T_2145 | _T_2139; // @[Mux.scala 27:72]
  wire  _T_2118 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2140 = _T_2118 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2147 = _T_2146 | _T_2140; // @[Mux.scala 27:72]
  wire  _T_2122 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2141 = _T_2122 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2148 = _T_2147 | _T_2141; // @[Mux.scala 27:72]
  wire  _T_2126 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2142 = _T_2126 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2149 = _T_2148 | _T_2142; // @[Mux.scala 27:72]
  wire  _T_2130 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2143 = _T_2130 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2150 = _T_2149 | _T_2143; // @[Mux.scala 27:72]
  wire  _T_2134 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2144 = _T_2134 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2150 | _T_2144; // @[Mux.scala 27:72]
  wire  _T_2192 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 453:69]
  wire  _T_2193 = ic_miss_buff_data_valid_bypass_index & _T_2192; // @[el2_ifu_mem_ctl.scala 453:67]
  wire  _T_2195 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 453:91]
  wire  _T_2196 = _T_2193 & _T_2195; // @[el2_ifu_mem_ctl.scala 453:89]
  wire  _T_2201 = _T_2193 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 454:65]
  wire  _T_2202 = _T_2196 | _T_2201; // @[el2_ifu_mem_ctl.scala 453:112]
  wire  _T_2204 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 455:43]
  wire  _T_2207 = _T_2204 & _T_2195; // @[el2_ifu_mem_ctl.scala 455:65]
  wire  _T_2208 = _T_2202 | _T_2207; // @[el2_ifu_mem_ctl.scala 454:88]
  wire  _T_2212 = _T_2204 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 456:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 433:75]
  wire  _T_2152 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2176 = _T_2152 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2155 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2177 = _T_2155 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2184 = _T_2176 | _T_2177; // @[Mux.scala 27:72]
  wire  _T_2158 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2178 = _T_2158 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2185 = _T_2184 | _T_2178; // @[Mux.scala 27:72]
  wire  _T_2161 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2179 = _T_2161 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2186 = _T_2185 | _T_2179; // @[Mux.scala 27:72]
  wire  _T_2164 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2180 = _T_2164 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2187 = _T_2186 | _T_2180; // @[Mux.scala 27:72]
  wire  _T_2167 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2181 = _T_2167 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2188 = _T_2187 | _T_2181; // @[Mux.scala 27:72]
  wire  _T_2170 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2182 = _T_2170 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2189 = _T_2188 | _T_2182; // @[Mux.scala 27:72]
  wire  _T_2173 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2183 = _T_2173 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2189 | _T_2183; // @[Mux.scala 27:72]
  wire  _T_2213 = _T_2212 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 456:87]
  wire  _T_2214 = _T_2208 | _T_2213; // @[el2_ifu_mem_ctl.scala 455:88]
  wire  _T_2218 = ic_miss_buff_data_valid_bypass_index & _T_2134; // @[el2_ifu_mem_ctl.scala 457:43]
  wire  miss_buff_hit_unq_f = _T_2214 | _T_2218; // @[el2_ifu_mem_ctl.scala 456:131]
  wire  _T_2234 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 462:55]
  wire  _T_2235 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 462:87]
  wire  _T_2236 = _T_2234 | _T_2235; // @[el2_ifu_mem_ctl.scala 462:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2236; // @[el2_ifu_mem_ctl.scala 462:41]
  wire  _T_2219 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 459:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 313:49]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[el2_ifu_mem_ctl.scala 450:51]
  wire  _T_2220 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 459:68]
  wire  _T_2221 = miss_buff_hit_unq_f & _T_2220; // @[el2_ifu_mem_ctl.scala 459:66]
  wire  stream_hit_f = _T_2219 & _T_2221; // @[el2_ifu_mem_ctl.scala 459:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 280:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 280:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 280:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 604:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 631:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 207:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 207:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 207:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 207:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 207:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 208:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 208:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 208:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 209:16]
  wire  _T_44 = _T_42 & _T_319; // @[el2_ifu_mem_ctl.scala 209:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 209:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 209:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 210:49]
  wire  _T_54 = ic_byp_hit_f & _T_319; // @[el2_ifu_mem_ctl.scala 211:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 211:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 211:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 199:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 211:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 211:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 211:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_319; // @[el2_ifu_mem_ctl.scala 212:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 212:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 212:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 212:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 213:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 214:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 214:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 214:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 213:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 212:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 211:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 210:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 209:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 208:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 207:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2231 = byp_fetch_index[4:1] == 4'hf; // @[el2_ifu_mem_ctl.scala 461:60]
  wire  _T_2232 = _T_2231 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 461:94]
  wire  stream_eol_f = _T_2232 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 461:112]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 222:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 222:87]
  wire  _T_113 = _T_111 & _T_2573; // @[el2_ifu_mem_ctl.scala 222:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 222:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 226:48]
  wire  _T_126 = _T_124 & _T_2573; // @[el2_ifu_mem_ctl.scala 226:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 226:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 286:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 286:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 286:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 286:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 286:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 287:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 286:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 287:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 341:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 287:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 287:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 287:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 230:50]
  wire  _T_137 = _T_135 & _T_2573; // @[el2_ifu_mem_ctl.scala 230:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 288:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 289:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 289:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 288:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 231:35]
  wire  _T_143 = _T_141 & _T_2573; // @[el2_ifu_mem_ctl.scala 231:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 231:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 230:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 236:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 235:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 235:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 240:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 240:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 197:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 197:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 197:26]
  wire  _T_30 = ic_act_miss_f & _T_2573; // @[el2_ifu_mem_ctl.scala 204:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 215:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 215:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 215:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 215:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 215:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 215:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 219:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 219:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 219:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 223:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 223:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 227:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 227:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 232:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 232:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 232:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 237:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 237:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 256:95]
  wire  _T_175 = _T_2234 & _T_174; // @[el2_ifu_mem_ctl.scala 256:93]
  wire  crit_wd_byp_ok_ff = _T_2235 | _T_175; // @[el2_ifu_mem_ctl.scala 256:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 257:36]
  wire  _T_180 = _T_2234 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 257:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 257:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 257:70]
  wire  _T_184 = _T_2234 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 258:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 258:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 257:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 258:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 259:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 259:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 258:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 261:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 261:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 269:64]
  reg [6:0] ifu_ic_rw_int_addr_ff; // @[el2_ifu_mem_ctl.scala 738:14]
  wire  _T_4619 = ifu_ic_rw_int_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_0; // @[Reg.scala 27:20]
  wire  _T_4747 = _T_4619 & way_status_out_0; // @[Mux.scala 27:72]
  wire  _T_4620 = ifu_ic_rw_int_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_1; // @[Reg.scala 27:20]
  wire  _T_4748 = _T_4620 & way_status_out_1; // @[Mux.scala 27:72]
  wire  _T_4875 = _T_4747 | _T_4748; // @[Mux.scala 27:72]
  wire  _T_4621 = ifu_ic_rw_int_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_2; // @[Reg.scala 27:20]
  wire  _T_4749 = _T_4621 & way_status_out_2; // @[Mux.scala 27:72]
  wire  _T_4876 = _T_4875 | _T_4749; // @[Mux.scala 27:72]
  wire  _T_4622 = ifu_ic_rw_int_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_3; // @[Reg.scala 27:20]
  wire  _T_4750 = _T_4622 & way_status_out_3; // @[Mux.scala 27:72]
  wire  _T_4877 = _T_4876 | _T_4750; // @[Mux.scala 27:72]
  wire  _T_4623 = ifu_ic_rw_int_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_4; // @[Reg.scala 27:20]
  wire  _T_4751 = _T_4623 & way_status_out_4; // @[Mux.scala 27:72]
  wire  _T_4878 = _T_4877 | _T_4751; // @[Mux.scala 27:72]
  wire  _T_4624 = ifu_ic_rw_int_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_5; // @[Reg.scala 27:20]
  wire  _T_4752 = _T_4624 & way_status_out_5; // @[Mux.scala 27:72]
  wire  _T_4879 = _T_4878 | _T_4752; // @[Mux.scala 27:72]
  wire  _T_4625 = ifu_ic_rw_int_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_6; // @[Reg.scala 27:20]
  wire  _T_4753 = _T_4625 & way_status_out_6; // @[Mux.scala 27:72]
  wire  _T_4880 = _T_4879 | _T_4753; // @[Mux.scala 27:72]
  wire  _T_4626 = ifu_ic_rw_int_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_7; // @[Reg.scala 27:20]
  wire  _T_4754 = _T_4626 & way_status_out_7; // @[Mux.scala 27:72]
  wire  _T_4881 = _T_4880 | _T_4754; // @[Mux.scala 27:72]
  wire  _T_4627 = ifu_ic_rw_int_addr_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_8; // @[Reg.scala 27:20]
  wire  _T_4755 = _T_4627 & way_status_out_8; // @[Mux.scala 27:72]
  wire  _T_4882 = _T_4881 | _T_4755; // @[Mux.scala 27:72]
  wire  _T_4628 = ifu_ic_rw_int_addr_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_9; // @[Reg.scala 27:20]
  wire  _T_4756 = _T_4628 & way_status_out_9; // @[Mux.scala 27:72]
  wire  _T_4883 = _T_4882 | _T_4756; // @[Mux.scala 27:72]
  wire  _T_4629 = ifu_ic_rw_int_addr_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_10; // @[Reg.scala 27:20]
  wire  _T_4757 = _T_4629 & way_status_out_10; // @[Mux.scala 27:72]
  wire  _T_4884 = _T_4883 | _T_4757; // @[Mux.scala 27:72]
  wire  _T_4630 = ifu_ic_rw_int_addr_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_11; // @[Reg.scala 27:20]
  wire  _T_4758 = _T_4630 & way_status_out_11; // @[Mux.scala 27:72]
  wire  _T_4885 = _T_4884 | _T_4758; // @[Mux.scala 27:72]
  wire  _T_4631 = ifu_ic_rw_int_addr_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_12; // @[Reg.scala 27:20]
  wire  _T_4759 = _T_4631 & way_status_out_12; // @[Mux.scala 27:72]
  wire  _T_4886 = _T_4885 | _T_4759; // @[Mux.scala 27:72]
  wire  _T_4632 = ifu_ic_rw_int_addr_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_13; // @[Reg.scala 27:20]
  wire  _T_4760 = _T_4632 & way_status_out_13; // @[Mux.scala 27:72]
  wire  _T_4887 = _T_4886 | _T_4760; // @[Mux.scala 27:72]
  wire  _T_4633 = ifu_ic_rw_int_addr_ff == 7'he; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_14; // @[Reg.scala 27:20]
  wire  _T_4761 = _T_4633 & way_status_out_14; // @[Mux.scala 27:72]
  wire  _T_4888 = _T_4887 | _T_4761; // @[Mux.scala 27:72]
  wire  _T_4634 = ifu_ic_rw_int_addr_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_15; // @[Reg.scala 27:20]
  wire  _T_4762 = _T_4634 & way_status_out_15; // @[Mux.scala 27:72]
  wire  _T_4889 = _T_4888 | _T_4762; // @[Mux.scala 27:72]
  wire  _T_4635 = ifu_ic_rw_int_addr_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_16; // @[Reg.scala 27:20]
  wire  _T_4763 = _T_4635 & way_status_out_16; // @[Mux.scala 27:72]
  wire  _T_4890 = _T_4889 | _T_4763; // @[Mux.scala 27:72]
  wire  _T_4636 = ifu_ic_rw_int_addr_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_17; // @[Reg.scala 27:20]
  wire  _T_4764 = _T_4636 & way_status_out_17; // @[Mux.scala 27:72]
  wire  _T_4891 = _T_4890 | _T_4764; // @[Mux.scala 27:72]
  wire  _T_4637 = ifu_ic_rw_int_addr_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_18; // @[Reg.scala 27:20]
  wire  _T_4765 = _T_4637 & way_status_out_18; // @[Mux.scala 27:72]
  wire  _T_4892 = _T_4891 | _T_4765; // @[Mux.scala 27:72]
  wire  _T_4638 = ifu_ic_rw_int_addr_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_19; // @[Reg.scala 27:20]
  wire  _T_4766 = _T_4638 & way_status_out_19; // @[Mux.scala 27:72]
  wire  _T_4893 = _T_4892 | _T_4766; // @[Mux.scala 27:72]
  wire  _T_4639 = ifu_ic_rw_int_addr_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_20; // @[Reg.scala 27:20]
  wire  _T_4767 = _T_4639 & way_status_out_20; // @[Mux.scala 27:72]
  wire  _T_4894 = _T_4893 | _T_4767; // @[Mux.scala 27:72]
  wire  _T_4640 = ifu_ic_rw_int_addr_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_21; // @[Reg.scala 27:20]
  wire  _T_4768 = _T_4640 & way_status_out_21; // @[Mux.scala 27:72]
  wire  _T_4895 = _T_4894 | _T_4768; // @[Mux.scala 27:72]
  wire  _T_4641 = ifu_ic_rw_int_addr_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_22; // @[Reg.scala 27:20]
  wire  _T_4769 = _T_4641 & way_status_out_22; // @[Mux.scala 27:72]
  wire  _T_4896 = _T_4895 | _T_4769; // @[Mux.scala 27:72]
  wire  _T_4642 = ifu_ic_rw_int_addr_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_23; // @[Reg.scala 27:20]
  wire  _T_4770 = _T_4642 & way_status_out_23; // @[Mux.scala 27:72]
  wire  _T_4897 = _T_4896 | _T_4770; // @[Mux.scala 27:72]
  wire  _T_4643 = ifu_ic_rw_int_addr_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_24; // @[Reg.scala 27:20]
  wire  _T_4771 = _T_4643 & way_status_out_24; // @[Mux.scala 27:72]
  wire  _T_4898 = _T_4897 | _T_4771; // @[Mux.scala 27:72]
  wire  _T_4644 = ifu_ic_rw_int_addr_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_25; // @[Reg.scala 27:20]
  wire  _T_4772 = _T_4644 & way_status_out_25; // @[Mux.scala 27:72]
  wire  _T_4899 = _T_4898 | _T_4772; // @[Mux.scala 27:72]
  wire  _T_4645 = ifu_ic_rw_int_addr_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_26; // @[Reg.scala 27:20]
  wire  _T_4773 = _T_4645 & way_status_out_26; // @[Mux.scala 27:72]
  wire  _T_4900 = _T_4899 | _T_4773; // @[Mux.scala 27:72]
  wire  _T_4646 = ifu_ic_rw_int_addr_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_27; // @[Reg.scala 27:20]
  wire  _T_4774 = _T_4646 & way_status_out_27; // @[Mux.scala 27:72]
  wire  _T_4901 = _T_4900 | _T_4774; // @[Mux.scala 27:72]
  wire  _T_4647 = ifu_ic_rw_int_addr_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_28; // @[Reg.scala 27:20]
  wire  _T_4775 = _T_4647 & way_status_out_28; // @[Mux.scala 27:72]
  wire  _T_4902 = _T_4901 | _T_4775; // @[Mux.scala 27:72]
  wire  _T_4648 = ifu_ic_rw_int_addr_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_29; // @[Reg.scala 27:20]
  wire  _T_4776 = _T_4648 & way_status_out_29; // @[Mux.scala 27:72]
  wire  _T_4903 = _T_4902 | _T_4776; // @[Mux.scala 27:72]
  wire  _T_4649 = ifu_ic_rw_int_addr_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_30; // @[Reg.scala 27:20]
  wire  _T_4777 = _T_4649 & way_status_out_30; // @[Mux.scala 27:72]
  wire  _T_4904 = _T_4903 | _T_4777; // @[Mux.scala 27:72]
  wire  _T_4650 = ifu_ic_rw_int_addr_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_31; // @[Reg.scala 27:20]
  wire  _T_4778 = _T_4650 & way_status_out_31; // @[Mux.scala 27:72]
  wire  _T_4905 = _T_4904 | _T_4778; // @[Mux.scala 27:72]
  wire  _T_4651 = ifu_ic_rw_int_addr_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_32; // @[Reg.scala 27:20]
  wire  _T_4779 = _T_4651 & way_status_out_32; // @[Mux.scala 27:72]
  wire  _T_4906 = _T_4905 | _T_4779; // @[Mux.scala 27:72]
  wire  _T_4652 = ifu_ic_rw_int_addr_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_33; // @[Reg.scala 27:20]
  wire  _T_4780 = _T_4652 & way_status_out_33; // @[Mux.scala 27:72]
  wire  _T_4907 = _T_4906 | _T_4780; // @[Mux.scala 27:72]
  wire  _T_4653 = ifu_ic_rw_int_addr_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_34; // @[Reg.scala 27:20]
  wire  _T_4781 = _T_4653 & way_status_out_34; // @[Mux.scala 27:72]
  wire  _T_4908 = _T_4907 | _T_4781; // @[Mux.scala 27:72]
  wire  _T_4654 = ifu_ic_rw_int_addr_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_35; // @[Reg.scala 27:20]
  wire  _T_4782 = _T_4654 & way_status_out_35; // @[Mux.scala 27:72]
  wire  _T_4909 = _T_4908 | _T_4782; // @[Mux.scala 27:72]
  wire  _T_4655 = ifu_ic_rw_int_addr_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_36; // @[Reg.scala 27:20]
  wire  _T_4783 = _T_4655 & way_status_out_36; // @[Mux.scala 27:72]
  wire  _T_4910 = _T_4909 | _T_4783; // @[Mux.scala 27:72]
  wire  _T_4656 = ifu_ic_rw_int_addr_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_37; // @[Reg.scala 27:20]
  wire  _T_4784 = _T_4656 & way_status_out_37; // @[Mux.scala 27:72]
  wire  _T_4911 = _T_4910 | _T_4784; // @[Mux.scala 27:72]
  wire  _T_4657 = ifu_ic_rw_int_addr_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_38; // @[Reg.scala 27:20]
  wire  _T_4785 = _T_4657 & way_status_out_38; // @[Mux.scala 27:72]
  wire  _T_4912 = _T_4911 | _T_4785; // @[Mux.scala 27:72]
  wire  _T_4658 = ifu_ic_rw_int_addr_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_39; // @[Reg.scala 27:20]
  wire  _T_4786 = _T_4658 & way_status_out_39; // @[Mux.scala 27:72]
  wire  _T_4913 = _T_4912 | _T_4786; // @[Mux.scala 27:72]
  wire  _T_4659 = ifu_ic_rw_int_addr_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_40; // @[Reg.scala 27:20]
  wire  _T_4787 = _T_4659 & way_status_out_40; // @[Mux.scala 27:72]
  wire  _T_4914 = _T_4913 | _T_4787; // @[Mux.scala 27:72]
  wire  _T_4660 = ifu_ic_rw_int_addr_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_41; // @[Reg.scala 27:20]
  wire  _T_4788 = _T_4660 & way_status_out_41; // @[Mux.scala 27:72]
  wire  _T_4915 = _T_4914 | _T_4788; // @[Mux.scala 27:72]
  wire  _T_4661 = ifu_ic_rw_int_addr_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_42; // @[Reg.scala 27:20]
  wire  _T_4789 = _T_4661 & way_status_out_42; // @[Mux.scala 27:72]
  wire  _T_4916 = _T_4915 | _T_4789; // @[Mux.scala 27:72]
  wire  _T_4662 = ifu_ic_rw_int_addr_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_43; // @[Reg.scala 27:20]
  wire  _T_4790 = _T_4662 & way_status_out_43; // @[Mux.scala 27:72]
  wire  _T_4917 = _T_4916 | _T_4790; // @[Mux.scala 27:72]
  wire  _T_4663 = ifu_ic_rw_int_addr_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_44; // @[Reg.scala 27:20]
  wire  _T_4791 = _T_4663 & way_status_out_44; // @[Mux.scala 27:72]
  wire  _T_4918 = _T_4917 | _T_4791; // @[Mux.scala 27:72]
  wire  _T_4664 = ifu_ic_rw_int_addr_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_45; // @[Reg.scala 27:20]
  wire  _T_4792 = _T_4664 & way_status_out_45; // @[Mux.scala 27:72]
  wire  _T_4919 = _T_4918 | _T_4792; // @[Mux.scala 27:72]
  wire  _T_4665 = ifu_ic_rw_int_addr_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_46; // @[Reg.scala 27:20]
  wire  _T_4793 = _T_4665 & way_status_out_46; // @[Mux.scala 27:72]
  wire  _T_4920 = _T_4919 | _T_4793; // @[Mux.scala 27:72]
  wire  _T_4666 = ifu_ic_rw_int_addr_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_47; // @[Reg.scala 27:20]
  wire  _T_4794 = _T_4666 & way_status_out_47; // @[Mux.scala 27:72]
  wire  _T_4921 = _T_4920 | _T_4794; // @[Mux.scala 27:72]
  wire  _T_4667 = ifu_ic_rw_int_addr_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_48; // @[Reg.scala 27:20]
  wire  _T_4795 = _T_4667 & way_status_out_48; // @[Mux.scala 27:72]
  wire  _T_4922 = _T_4921 | _T_4795; // @[Mux.scala 27:72]
  wire  _T_4668 = ifu_ic_rw_int_addr_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_49; // @[Reg.scala 27:20]
  wire  _T_4796 = _T_4668 & way_status_out_49; // @[Mux.scala 27:72]
  wire  _T_4923 = _T_4922 | _T_4796; // @[Mux.scala 27:72]
  wire  _T_4669 = ifu_ic_rw_int_addr_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_50; // @[Reg.scala 27:20]
  wire  _T_4797 = _T_4669 & way_status_out_50; // @[Mux.scala 27:72]
  wire  _T_4924 = _T_4923 | _T_4797; // @[Mux.scala 27:72]
  wire  _T_4670 = ifu_ic_rw_int_addr_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_51; // @[Reg.scala 27:20]
  wire  _T_4798 = _T_4670 & way_status_out_51; // @[Mux.scala 27:72]
  wire  _T_4925 = _T_4924 | _T_4798; // @[Mux.scala 27:72]
  wire  _T_4671 = ifu_ic_rw_int_addr_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_52; // @[Reg.scala 27:20]
  wire  _T_4799 = _T_4671 & way_status_out_52; // @[Mux.scala 27:72]
  wire  _T_4926 = _T_4925 | _T_4799; // @[Mux.scala 27:72]
  wire  _T_4672 = ifu_ic_rw_int_addr_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_53; // @[Reg.scala 27:20]
  wire  _T_4800 = _T_4672 & way_status_out_53; // @[Mux.scala 27:72]
  wire  _T_4927 = _T_4926 | _T_4800; // @[Mux.scala 27:72]
  wire  _T_4673 = ifu_ic_rw_int_addr_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_54; // @[Reg.scala 27:20]
  wire  _T_4801 = _T_4673 & way_status_out_54; // @[Mux.scala 27:72]
  wire  _T_4928 = _T_4927 | _T_4801; // @[Mux.scala 27:72]
  wire  _T_4674 = ifu_ic_rw_int_addr_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_55; // @[Reg.scala 27:20]
  wire  _T_4802 = _T_4674 & way_status_out_55; // @[Mux.scala 27:72]
  wire  _T_4929 = _T_4928 | _T_4802; // @[Mux.scala 27:72]
  wire  _T_4675 = ifu_ic_rw_int_addr_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_56; // @[Reg.scala 27:20]
  wire  _T_4803 = _T_4675 & way_status_out_56; // @[Mux.scala 27:72]
  wire  _T_4930 = _T_4929 | _T_4803; // @[Mux.scala 27:72]
  wire  _T_4676 = ifu_ic_rw_int_addr_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_57; // @[Reg.scala 27:20]
  wire  _T_4804 = _T_4676 & way_status_out_57; // @[Mux.scala 27:72]
  wire  _T_4931 = _T_4930 | _T_4804; // @[Mux.scala 27:72]
  wire  _T_4677 = ifu_ic_rw_int_addr_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_58; // @[Reg.scala 27:20]
  wire  _T_4805 = _T_4677 & way_status_out_58; // @[Mux.scala 27:72]
  wire  _T_4932 = _T_4931 | _T_4805; // @[Mux.scala 27:72]
  wire  _T_4678 = ifu_ic_rw_int_addr_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_59; // @[Reg.scala 27:20]
  wire  _T_4806 = _T_4678 & way_status_out_59; // @[Mux.scala 27:72]
  wire  _T_4933 = _T_4932 | _T_4806; // @[Mux.scala 27:72]
  wire  _T_4679 = ifu_ic_rw_int_addr_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_60; // @[Reg.scala 27:20]
  wire  _T_4807 = _T_4679 & way_status_out_60; // @[Mux.scala 27:72]
  wire  _T_4934 = _T_4933 | _T_4807; // @[Mux.scala 27:72]
  wire  _T_4680 = ifu_ic_rw_int_addr_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_61; // @[Reg.scala 27:20]
  wire  _T_4808 = _T_4680 & way_status_out_61; // @[Mux.scala 27:72]
  wire  _T_4935 = _T_4934 | _T_4808; // @[Mux.scala 27:72]
  wire  _T_4681 = ifu_ic_rw_int_addr_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_62; // @[Reg.scala 27:20]
  wire  _T_4809 = _T_4681 & way_status_out_62; // @[Mux.scala 27:72]
  wire  _T_4936 = _T_4935 | _T_4809; // @[Mux.scala 27:72]
  wire  _T_4682 = ifu_ic_rw_int_addr_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_63; // @[Reg.scala 27:20]
  wire  _T_4810 = _T_4682 & way_status_out_63; // @[Mux.scala 27:72]
  wire  _T_4937 = _T_4936 | _T_4810; // @[Mux.scala 27:72]
  wire  _T_4683 = ifu_ic_rw_int_addr_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_64; // @[Reg.scala 27:20]
  wire  _T_4811 = _T_4683 & way_status_out_64; // @[Mux.scala 27:72]
  wire  _T_4938 = _T_4937 | _T_4811; // @[Mux.scala 27:72]
  wire  _T_4684 = ifu_ic_rw_int_addr_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_65; // @[Reg.scala 27:20]
  wire  _T_4812 = _T_4684 & way_status_out_65; // @[Mux.scala 27:72]
  wire  _T_4939 = _T_4938 | _T_4812; // @[Mux.scala 27:72]
  wire  _T_4685 = ifu_ic_rw_int_addr_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_66; // @[Reg.scala 27:20]
  wire  _T_4813 = _T_4685 & way_status_out_66; // @[Mux.scala 27:72]
  wire  _T_4940 = _T_4939 | _T_4813; // @[Mux.scala 27:72]
  wire  _T_4686 = ifu_ic_rw_int_addr_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_67; // @[Reg.scala 27:20]
  wire  _T_4814 = _T_4686 & way_status_out_67; // @[Mux.scala 27:72]
  wire  _T_4941 = _T_4940 | _T_4814; // @[Mux.scala 27:72]
  wire  _T_4687 = ifu_ic_rw_int_addr_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_68; // @[Reg.scala 27:20]
  wire  _T_4815 = _T_4687 & way_status_out_68; // @[Mux.scala 27:72]
  wire  _T_4942 = _T_4941 | _T_4815; // @[Mux.scala 27:72]
  wire  _T_4688 = ifu_ic_rw_int_addr_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_69; // @[Reg.scala 27:20]
  wire  _T_4816 = _T_4688 & way_status_out_69; // @[Mux.scala 27:72]
  wire  _T_4943 = _T_4942 | _T_4816; // @[Mux.scala 27:72]
  wire  _T_4689 = ifu_ic_rw_int_addr_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_70; // @[Reg.scala 27:20]
  wire  _T_4817 = _T_4689 & way_status_out_70; // @[Mux.scala 27:72]
  wire  _T_4944 = _T_4943 | _T_4817; // @[Mux.scala 27:72]
  wire  _T_4690 = ifu_ic_rw_int_addr_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_71; // @[Reg.scala 27:20]
  wire  _T_4818 = _T_4690 & way_status_out_71; // @[Mux.scala 27:72]
  wire  _T_4945 = _T_4944 | _T_4818; // @[Mux.scala 27:72]
  wire  _T_4691 = ifu_ic_rw_int_addr_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_72; // @[Reg.scala 27:20]
  wire  _T_4819 = _T_4691 & way_status_out_72; // @[Mux.scala 27:72]
  wire  _T_4946 = _T_4945 | _T_4819; // @[Mux.scala 27:72]
  wire  _T_4692 = ifu_ic_rw_int_addr_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_73; // @[Reg.scala 27:20]
  wire  _T_4820 = _T_4692 & way_status_out_73; // @[Mux.scala 27:72]
  wire  _T_4947 = _T_4946 | _T_4820; // @[Mux.scala 27:72]
  wire  _T_4693 = ifu_ic_rw_int_addr_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_74; // @[Reg.scala 27:20]
  wire  _T_4821 = _T_4693 & way_status_out_74; // @[Mux.scala 27:72]
  wire  _T_4948 = _T_4947 | _T_4821; // @[Mux.scala 27:72]
  wire  _T_4694 = ifu_ic_rw_int_addr_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_75; // @[Reg.scala 27:20]
  wire  _T_4822 = _T_4694 & way_status_out_75; // @[Mux.scala 27:72]
  wire  _T_4949 = _T_4948 | _T_4822; // @[Mux.scala 27:72]
  wire  _T_4695 = ifu_ic_rw_int_addr_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_76; // @[Reg.scala 27:20]
  wire  _T_4823 = _T_4695 & way_status_out_76; // @[Mux.scala 27:72]
  wire  _T_4950 = _T_4949 | _T_4823; // @[Mux.scala 27:72]
  wire  _T_4696 = ifu_ic_rw_int_addr_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_77; // @[Reg.scala 27:20]
  wire  _T_4824 = _T_4696 & way_status_out_77; // @[Mux.scala 27:72]
  wire  _T_4951 = _T_4950 | _T_4824; // @[Mux.scala 27:72]
  wire  _T_4697 = ifu_ic_rw_int_addr_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_78; // @[Reg.scala 27:20]
  wire  _T_4825 = _T_4697 & way_status_out_78; // @[Mux.scala 27:72]
  wire  _T_4952 = _T_4951 | _T_4825; // @[Mux.scala 27:72]
  wire  _T_4698 = ifu_ic_rw_int_addr_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_79; // @[Reg.scala 27:20]
  wire  _T_4826 = _T_4698 & way_status_out_79; // @[Mux.scala 27:72]
  wire  _T_4953 = _T_4952 | _T_4826; // @[Mux.scala 27:72]
  wire  _T_4699 = ifu_ic_rw_int_addr_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_80; // @[Reg.scala 27:20]
  wire  _T_4827 = _T_4699 & way_status_out_80; // @[Mux.scala 27:72]
  wire  _T_4954 = _T_4953 | _T_4827; // @[Mux.scala 27:72]
  wire  _T_4700 = ifu_ic_rw_int_addr_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_81; // @[Reg.scala 27:20]
  wire  _T_4828 = _T_4700 & way_status_out_81; // @[Mux.scala 27:72]
  wire  _T_4955 = _T_4954 | _T_4828; // @[Mux.scala 27:72]
  wire  _T_4701 = ifu_ic_rw_int_addr_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_82; // @[Reg.scala 27:20]
  wire  _T_4829 = _T_4701 & way_status_out_82; // @[Mux.scala 27:72]
  wire  _T_4956 = _T_4955 | _T_4829; // @[Mux.scala 27:72]
  wire  _T_4702 = ifu_ic_rw_int_addr_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_83; // @[Reg.scala 27:20]
  wire  _T_4830 = _T_4702 & way_status_out_83; // @[Mux.scala 27:72]
  wire  _T_4957 = _T_4956 | _T_4830; // @[Mux.scala 27:72]
  wire  _T_4703 = ifu_ic_rw_int_addr_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_84; // @[Reg.scala 27:20]
  wire  _T_4831 = _T_4703 & way_status_out_84; // @[Mux.scala 27:72]
  wire  _T_4958 = _T_4957 | _T_4831; // @[Mux.scala 27:72]
  wire  _T_4704 = ifu_ic_rw_int_addr_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_85; // @[Reg.scala 27:20]
  wire  _T_4832 = _T_4704 & way_status_out_85; // @[Mux.scala 27:72]
  wire  _T_4959 = _T_4958 | _T_4832; // @[Mux.scala 27:72]
  wire  _T_4705 = ifu_ic_rw_int_addr_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_86; // @[Reg.scala 27:20]
  wire  _T_4833 = _T_4705 & way_status_out_86; // @[Mux.scala 27:72]
  wire  _T_4960 = _T_4959 | _T_4833; // @[Mux.scala 27:72]
  wire  _T_4706 = ifu_ic_rw_int_addr_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_87; // @[Reg.scala 27:20]
  wire  _T_4834 = _T_4706 & way_status_out_87; // @[Mux.scala 27:72]
  wire  _T_4961 = _T_4960 | _T_4834; // @[Mux.scala 27:72]
  wire  _T_4707 = ifu_ic_rw_int_addr_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_88; // @[Reg.scala 27:20]
  wire  _T_4835 = _T_4707 & way_status_out_88; // @[Mux.scala 27:72]
  wire  _T_4962 = _T_4961 | _T_4835; // @[Mux.scala 27:72]
  wire  _T_4708 = ifu_ic_rw_int_addr_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_89; // @[Reg.scala 27:20]
  wire  _T_4836 = _T_4708 & way_status_out_89; // @[Mux.scala 27:72]
  wire  _T_4963 = _T_4962 | _T_4836; // @[Mux.scala 27:72]
  wire  _T_4709 = ifu_ic_rw_int_addr_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_90; // @[Reg.scala 27:20]
  wire  _T_4837 = _T_4709 & way_status_out_90; // @[Mux.scala 27:72]
  wire  _T_4964 = _T_4963 | _T_4837; // @[Mux.scala 27:72]
  wire  _T_4710 = ifu_ic_rw_int_addr_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_91; // @[Reg.scala 27:20]
  wire  _T_4838 = _T_4710 & way_status_out_91; // @[Mux.scala 27:72]
  wire  _T_4965 = _T_4964 | _T_4838; // @[Mux.scala 27:72]
  wire  _T_4711 = ifu_ic_rw_int_addr_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_92; // @[Reg.scala 27:20]
  wire  _T_4839 = _T_4711 & way_status_out_92; // @[Mux.scala 27:72]
  wire  _T_4966 = _T_4965 | _T_4839; // @[Mux.scala 27:72]
  wire  _T_4712 = ifu_ic_rw_int_addr_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_93; // @[Reg.scala 27:20]
  wire  _T_4840 = _T_4712 & way_status_out_93; // @[Mux.scala 27:72]
  wire  _T_4967 = _T_4966 | _T_4840; // @[Mux.scala 27:72]
  wire  _T_4713 = ifu_ic_rw_int_addr_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_94; // @[Reg.scala 27:20]
  wire  _T_4841 = _T_4713 & way_status_out_94; // @[Mux.scala 27:72]
  wire  _T_4968 = _T_4967 | _T_4841; // @[Mux.scala 27:72]
  wire  _T_4714 = ifu_ic_rw_int_addr_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_95; // @[Reg.scala 27:20]
  wire  _T_4842 = _T_4714 & way_status_out_95; // @[Mux.scala 27:72]
  wire  _T_4969 = _T_4968 | _T_4842; // @[Mux.scala 27:72]
  wire  _T_4715 = ifu_ic_rw_int_addr_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_96; // @[Reg.scala 27:20]
  wire  _T_4843 = _T_4715 & way_status_out_96; // @[Mux.scala 27:72]
  wire  _T_4970 = _T_4969 | _T_4843; // @[Mux.scala 27:72]
  wire  _T_4716 = ifu_ic_rw_int_addr_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_97; // @[Reg.scala 27:20]
  wire  _T_4844 = _T_4716 & way_status_out_97; // @[Mux.scala 27:72]
  wire  _T_4971 = _T_4970 | _T_4844; // @[Mux.scala 27:72]
  wire  _T_4717 = ifu_ic_rw_int_addr_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_98; // @[Reg.scala 27:20]
  wire  _T_4845 = _T_4717 & way_status_out_98; // @[Mux.scala 27:72]
  wire  _T_4972 = _T_4971 | _T_4845; // @[Mux.scala 27:72]
  wire  _T_4718 = ifu_ic_rw_int_addr_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_99; // @[Reg.scala 27:20]
  wire  _T_4846 = _T_4718 & way_status_out_99; // @[Mux.scala 27:72]
  wire  _T_4973 = _T_4972 | _T_4846; // @[Mux.scala 27:72]
  wire  _T_4719 = ifu_ic_rw_int_addr_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_100; // @[Reg.scala 27:20]
  wire  _T_4847 = _T_4719 & way_status_out_100; // @[Mux.scala 27:72]
  wire  _T_4974 = _T_4973 | _T_4847; // @[Mux.scala 27:72]
  wire  _T_4720 = ifu_ic_rw_int_addr_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_101; // @[Reg.scala 27:20]
  wire  _T_4848 = _T_4720 & way_status_out_101; // @[Mux.scala 27:72]
  wire  _T_4975 = _T_4974 | _T_4848; // @[Mux.scala 27:72]
  wire  _T_4721 = ifu_ic_rw_int_addr_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_102; // @[Reg.scala 27:20]
  wire  _T_4849 = _T_4721 & way_status_out_102; // @[Mux.scala 27:72]
  wire  _T_4976 = _T_4975 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4722 = ifu_ic_rw_int_addr_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_103; // @[Reg.scala 27:20]
  wire  _T_4850 = _T_4722 & way_status_out_103; // @[Mux.scala 27:72]
  wire  _T_4977 = _T_4976 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4723 = ifu_ic_rw_int_addr_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_104; // @[Reg.scala 27:20]
  wire  _T_4851 = _T_4723 & way_status_out_104; // @[Mux.scala 27:72]
  wire  _T_4978 = _T_4977 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_4724 = ifu_ic_rw_int_addr_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_105; // @[Reg.scala 27:20]
  wire  _T_4852 = _T_4724 & way_status_out_105; // @[Mux.scala 27:72]
  wire  _T_4979 = _T_4978 | _T_4852; // @[Mux.scala 27:72]
  wire  _T_4725 = ifu_ic_rw_int_addr_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_106; // @[Reg.scala 27:20]
  wire  _T_4853 = _T_4725 & way_status_out_106; // @[Mux.scala 27:72]
  wire  _T_4980 = _T_4979 | _T_4853; // @[Mux.scala 27:72]
  wire  _T_4726 = ifu_ic_rw_int_addr_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_107; // @[Reg.scala 27:20]
  wire  _T_4854 = _T_4726 & way_status_out_107; // @[Mux.scala 27:72]
  wire  _T_4981 = _T_4980 | _T_4854; // @[Mux.scala 27:72]
  wire  _T_4727 = ifu_ic_rw_int_addr_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_108; // @[Reg.scala 27:20]
  wire  _T_4855 = _T_4727 & way_status_out_108; // @[Mux.scala 27:72]
  wire  _T_4982 = _T_4981 | _T_4855; // @[Mux.scala 27:72]
  wire  _T_4728 = ifu_ic_rw_int_addr_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_109; // @[Reg.scala 27:20]
  wire  _T_4856 = _T_4728 & way_status_out_109; // @[Mux.scala 27:72]
  wire  _T_4983 = _T_4982 | _T_4856; // @[Mux.scala 27:72]
  wire  _T_4729 = ifu_ic_rw_int_addr_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_110; // @[Reg.scala 27:20]
  wire  _T_4857 = _T_4729 & way_status_out_110; // @[Mux.scala 27:72]
  wire  _T_4984 = _T_4983 | _T_4857; // @[Mux.scala 27:72]
  wire  _T_4730 = ifu_ic_rw_int_addr_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_111; // @[Reg.scala 27:20]
  wire  _T_4858 = _T_4730 & way_status_out_111; // @[Mux.scala 27:72]
  wire  _T_4985 = _T_4984 | _T_4858; // @[Mux.scala 27:72]
  wire  _T_4731 = ifu_ic_rw_int_addr_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_112; // @[Reg.scala 27:20]
  wire  _T_4859 = _T_4731 & way_status_out_112; // @[Mux.scala 27:72]
  wire  _T_4986 = _T_4985 | _T_4859; // @[Mux.scala 27:72]
  wire  _T_4732 = ifu_ic_rw_int_addr_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_113; // @[Reg.scala 27:20]
  wire  _T_4860 = _T_4732 & way_status_out_113; // @[Mux.scala 27:72]
  wire  _T_4987 = _T_4986 | _T_4860; // @[Mux.scala 27:72]
  wire  _T_4733 = ifu_ic_rw_int_addr_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_114; // @[Reg.scala 27:20]
  wire  _T_4861 = _T_4733 & way_status_out_114; // @[Mux.scala 27:72]
  wire  _T_4988 = _T_4987 | _T_4861; // @[Mux.scala 27:72]
  wire  _T_4734 = ifu_ic_rw_int_addr_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_115; // @[Reg.scala 27:20]
  wire  _T_4862 = _T_4734 & way_status_out_115; // @[Mux.scala 27:72]
  wire  _T_4989 = _T_4988 | _T_4862; // @[Mux.scala 27:72]
  wire  _T_4735 = ifu_ic_rw_int_addr_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_116; // @[Reg.scala 27:20]
  wire  _T_4863 = _T_4735 & way_status_out_116; // @[Mux.scala 27:72]
  wire  _T_4990 = _T_4989 | _T_4863; // @[Mux.scala 27:72]
  wire  _T_4736 = ifu_ic_rw_int_addr_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_117; // @[Reg.scala 27:20]
  wire  _T_4864 = _T_4736 & way_status_out_117; // @[Mux.scala 27:72]
  wire  _T_4991 = _T_4990 | _T_4864; // @[Mux.scala 27:72]
  wire  _T_4737 = ifu_ic_rw_int_addr_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_118; // @[Reg.scala 27:20]
  wire  _T_4865 = _T_4737 & way_status_out_118; // @[Mux.scala 27:72]
  wire  _T_4992 = _T_4991 | _T_4865; // @[Mux.scala 27:72]
  wire  _T_4738 = ifu_ic_rw_int_addr_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_119; // @[Reg.scala 27:20]
  wire  _T_4866 = _T_4738 & way_status_out_119; // @[Mux.scala 27:72]
  wire  _T_4993 = _T_4992 | _T_4866; // @[Mux.scala 27:72]
  wire  _T_4739 = ifu_ic_rw_int_addr_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_120; // @[Reg.scala 27:20]
  wire  _T_4867 = _T_4739 & way_status_out_120; // @[Mux.scala 27:72]
  wire  _T_4994 = _T_4993 | _T_4867; // @[Mux.scala 27:72]
  wire  _T_4740 = ifu_ic_rw_int_addr_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_121; // @[Reg.scala 27:20]
  wire  _T_4868 = _T_4740 & way_status_out_121; // @[Mux.scala 27:72]
  wire  _T_4995 = _T_4994 | _T_4868; // @[Mux.scala 27:72]
  wire  _T_4741 = ifu_ic_rw_int_addr_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_122; // @[Reg.scala 27:20]
  wire  _T_4869 = _T_4741 & way_status_out_122; // @[Mux.scala 27:72]
  wire  _T_4996 = _T_4995 | _T_4869; // @[Mux.scala 27:72]
  wire  _T_4742 = ifu_ic_rw_int_addr_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_123; // @[Reg.scala 27:20]
  wire  _T_4870 = _T_4742 & way_status_out_123; // @[Mux.scala 27:72]
  wire  _T_4997 = _T_4996 | _T_4870; // @[Mux.scala 27:72]
  wire  _T_4743 = ifu_ic_rw_int_addr_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_124; // @[Reg.scala 27:20]
  wire  _T_4871 = _T_4743 & way_status_out_124; // @[Mux.scala 27:72]
  wire  _T_4998 = _T_4997 | _T_4871; // @[Mux.scala 27:72]
  wire  _T_4744 = ifu_ic_rw_int_addr_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_125; // @[Reg.scala 27:20]
  wire  _T_4872 = _T_4744 & way_status_out_125; // @[Mux.scala 27:72]
  wire  _T_4999 = _T_4998 | _T_4872; // @[Mux.scala 27:72]
  wire  _T_4745 = ifu_ic_rw_int_addr_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_126; // @[Reg.scala 27:20]
  wire  _T_4873 = _T_4745 & way_status_out_126; // @[Mux.scala 27:72]
  wire  _T_5000 = _T_4999 | _T_4873; // @[Mux.scala 27:72]
  wire  _T_4746 = ifu_ic_rw_int_addr_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 734:80]
  reg  way_status_out_127; // @[Reg.scala 27:20]
  wire  _T_4874 = _T_4746 & way_status_out_127; // @[Mux.scala 27:72]
  wire  way_status = _T_5000 | _T_4874; // @[Mux.scala 27:72]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 264:96]
  wire [1:0] _T_197 = _T_195 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_198 = _T_197 & io_ic_tag_valid; // @[el2_ifu_mem_ctl.scala 264:113]
  reg [1:0] tagv_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 270:58]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 266:67]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:54]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[el2_ifu_mem_ctl.scala 584:46]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 273:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 278:59]
  wire  _T_214 = _T_212 | _T_2219; // @[el2_ifu_mem_ctl.scala 278:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 278:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 284:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 284:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 284:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 284:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 291:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 291:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 291:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 292:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 292:32]
  wire  _T_274 = imb_ff[11:5] == imb_scnd_ff[11:5]; // @[el2_ifu_mem_ctl.scala 295:79]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 295:135]
  reg [1:0] ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 582:51]
  wire  _T_2643 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 627:48]
  wire  _T_2644 = _T_2643 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 627:52]
  wire  bus_ifu_wr_data_error_ff = _T_2644 & miss_pending; // @[el2_ifu_mem_ctl.scala 627:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 369:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 368:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 295:153]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 295:151]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 298:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 298:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 299:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 319:59]
  wire  _T_9704 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 790:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 320:53]
  wire  _T_9706 = _T_9704 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 790:51]
  wire  _T_9708 = _T_9706 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 790:67]
  wire  _T_9710 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 790:86]
  wire  replace_way_mb_any_0 = _T_9708 | _T_9710; // @[el2_ifu_mem_ctl.scala 790:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9713 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 791:50]
  wire  _T_9715 = _T_9713 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 791:66]
  wire  _T_9717 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 791:85]
  wire  _T_9719 = _T_9717 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 791:100]
  wire  replace_way_mb_any_1 = _T_9715 | _T_9719; // @[el2_ifu_mem_ctl.scala 791:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 303:110]
  wire [1:0] _T_290 = tagv_mb_scnd_ff | _T_289; // @[el2_ifu_mem_ctl.scala 303:62]
  wire [1:0] _T_295 = io_ic_tag_valid & _T_197; // @[el2_ifu_mem_ctl.scala 304:56]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 307:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 307:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 308:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 307:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 307:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 309:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 318:48]
  wire  _T_309 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 317:57]
  wire  _T_315 = _T_2234 & flush_final_f; // @[el2_ifu_mem_ctl.scala 322:87]
  wire  _T_316 = ~_T_315; // @[el2_ifu_mem_ctl.scala 322:55]
  wire  _T_317 = io_ifc_fetch_req_bf & _T_316; // @[el2_ifu_mem_ctl.scala 322:53]
  wire  _T_2226 = ~_T_2221; // @[el2_ifu_mem_ctl.scala 460:46]
  wire  _T_2227 = _T_2219 & _T_2226; // @[el2_ifu_mem_ctl.scala 460:44]
  wire  stream_miss_f = _T_2227 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 460:84]
  wire  _T_318 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 322:106]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 328:68]
  reg [2:0] bus_rd_addr_count; // @[el2_ifu_mem_ctl.scala 609:55]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_325 = _T_239 | _T_2219; // @[el2_ifu_mem_ctl.scala 330:55]
  wire  _T_328 = _T_325 & _T_56; // @[el2_ifu_mem_ctl.scala 330:82]
  wire  _T_2240 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 465:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2240}; // @[Cat.scala 29:58]
  wire  _T_2241 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2265 = _T_2241 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2244 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2266 = _T_2244 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2273 = _T_2265 | _T_2266; // @[Mux.scala 27:72]
  wire  _T_2247 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2267 = _T_2247 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2274 = _T_2273 | _T_2267; // @[Mux.scala 27:72]
  wire  _T_2250 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2268 = _T_2250 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2275 = _T_2274 | _T_2268; // @[Mux.scala 27:72]
  wire  _T_2253 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2269 = _T_2253 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2276 = _T_2275 | _T_2269; // @[Mux.scala 27:72]
  wire  _T_2256 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2270 = _T_2256 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2277 = _T_2276 | _T_2270; // @[Mux.scala 27:72]
  wire  _T_2259 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2271 = _T_2259 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2278 = _T_2277 | _T_2271; // @[Mux.scala 27:72]
  wire  _T_2262 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2272 = _T_2262 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2278 | _T_2272; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 467:46]
  wire  _T_332 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 334:35]
  wire  _T_334 = _T_332 & _T_17; // @[el2_ifu_mem_ctl.scala 334:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 624:61]
  wire  _T_2637 = ic_act_miss_f_delayed & _T_2235; // @[el2_ifu_mem_ctl.scala 625:53]
  wire  reset_tag_valid_for_miss = _T_2637 & _T_17; // @[el2_ifu_mem_ctl.scala 625:84]
  wire  sel_mb_addr = _T_334 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 334:79]
  wire [30:0] _T_338 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_339 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 336:37]
  wire [30:0] _T_340 = sel_mb_addr ? _T_338 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_341 = _T_339 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_340 | _T_341; // @[Mux.scala 27:72]
  wire  _T_346 = _T_334 & last_beat; // @[el2_ifu_mem_ctl.scala 338:84]
  wire  _T_2631 = ~_T_2643; // @[el2_ifu_mem_ctl.scala 622:84]
  wire  _T_2632 = _T_100 & _T_2631; // @[el2_ifu_mem_ctl.scala 622:82]
  wire  bus_ifu_wr_en_ff_q = _T_2632 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 622:108]
  wire  sel_mb_status_addr = _T_346 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 338:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_338 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 339:31]
  reg [63:0] ifu_bus_rdata_ff; // @[el2_ifu_mem_ctl.scala 583:48]
  wire [6:0] _T_569 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 416:13]
  wire  _T_570 = ^_T_569; // @[el2_lib.scala 416:20]
  wire [6:0] _T_576 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_583 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 416:30]
  wire [14:0] _T_584 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_576}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_591 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 416:30]
  wire [30:0] _T_600 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_591,_T_584}; // @[el2_lib.scala 416:30]
  wire  _T_601 = ^_T_600; // @[el2_lib.scala 416:37]
  wire [6:0] _T_607 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 416:47]
  wire [14:0] _T_615 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_607}; // @[el2_lib.scala 416:47]
  wire [30:0] _T_631 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_591,_T_615}; // @[el2_lib.scala 416:47]
  wire  _T_632 = ^_T_631; // @[el2_lib.scala 416:54]
  wire [6:0] _T_638 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 416:64]
  wire [14:0] _T_646 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_638}; // @[el2_lib.scala 416:64]
  wire [30:0] _T_662 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_583,_T_646}; // @[el2_lib.scala 416:64]
  wire  _T_663 = ^_T_662; // @[el2_lib.scala 416:71]
  wire [7:0] _T_670 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 416:81]
  wire [16:0] _T_679 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_670}; // @[el2_lib.scala 416:81]
  wire [8:0] _T_687 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 416:81]
  wire [17:0] _T_696 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_687}; // @[el2_lib.scala 416:81]
  wire [34:0] _T_697 = {_T_696,_T_679}; // @[el2_lib.scala 416:81]
  wire  _T_698 = ^_T_697; // @[el2_lib.scala 416:88]
  wire [7:0] _T_705 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 416:98]
  wire [16:0] _T_714 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_705}; // @[el2_lib.scala 416:98]
  wire [8:0] _T_722 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 416:98]
  wire [17:0] _T_731 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_722}; // @[el2_lib.scala 416:98]
  wire [34:0] _T_732 = {_T_731,_T_714}; // @[el2_lib.scala 416:98]
  wire  _T_733 = ^_T_732; // @[el2_lib.scala 416:105]
  wire [7:0] _T_740 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 416:115]
  wire [16:0] _T_749 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_740}; // @[el2_lib.scala 416:115]
  wire [8:0] _T_757 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 416:115]
  wire [17:0] _T_766 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_757}; // @[el2_lib.scala 416:115]
  wire [34:0] _T_767 = {_T_766,_T_749}; // @[el2_lib.scala 416:115]
  wire  _T_768 = ^_T_767; // @[el2_lib.scala 416:122]
  wire [3:0] _T_2281 = {ifu_bus_rid_ff[2:1],_T_2240,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2282 = _T_2281 == 4'h0; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_0; // @[el2_ifu_mem_ctl.scala 403:65]
  wire [31:0] _T_2329 = _T_2282 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2285 = _T_2281 == 4'h1; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_1; // @[el2_ifu_mem_ctl.scala 404:67]
  wire [31:0] _T_2330 = _T_2285 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2345 = _T_2329 | _T_2330; // @[Mux.scala 27:72]
  wire  _T_2288 = _T_2281 == 4'h2; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_2; // @[el2_ifu_mem_ctl.scala 403:65]
  wire [31:0] _T_2331 = _T_2288 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2346 = _T_2345 | _T_2331; // @[Mux.scala 27:72]
  wire  _T_2291 = _T_2281 == 4'h3; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_3; // @[el2_ifu_mem_ctl.scala 404:67]
  wire [31:0] _T_2332 = _T_2291 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2347 = _T_2346 | _T_2332; // @[Mux.scala 27:72]
  wire  _T_2294 = _T_2281 == 4'h4; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_4; // @[el2_ifu_mem_ctl.scala 403:65]
  wire [31:0] _T_2333 = _T_2294 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2348 = _T_2347 | _T_2333; // @[Mux.scala 27:72]
  wire  _T_2297 = _T_2281 == 4'h5; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_5; // @[el2_ifu_mem_ctl.scala 404:67]
  wire [31:0] _T_2334 = _T_2297 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2349 = _T_2348 | _T_2334; // @[Mux.scala 27:72]
  wire  _T_2300 = _T_2281 == 4'h6; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_6; // @[el2_ifu_mem_ctl.scala 403:65]
  wire [31:0] _T_2335 = _T_2300 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2350 = _T_2349 | _T_2335; // @[Mux.scala 27:72]
  wire  _T_2303 = _T_2281 == 4'h7; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_7; // @[el2_ifu_mem_ctl.scala 404:67]
  wire [31:0] _T_2336 = _T_2303 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2351 = _T_2350 | _T_2336; // @[Mux.scala 27:72]
  wire  _T_2306 = _T_2281 == 4'h8; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_8; // @[el2_ifu_mem_ctl.scala 403:65]
  wire [31:0] _T_2337 = _T_2306 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2352 = _T_2351 | _T_2337; // @[Mux.scala 27:72]
  wire  _T_2309 = _T_2281 == 4'h9; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_9; // @[el2_ifu_mem_ctl.scala 404:67]
  wire [31:0] _T_2338 = _T_2309 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2353 = _T_2352 | _T_2338; // @[Mux.scala 27:72]
  wire  _T_2312 = _T_2281 == 4'ha; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_10; // @[el2_ifu_mem_ctl.scala 403:65]
  wire [31:0] _T_2339 = _T_2312 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2354 = _T_2353 | _T_2339; // @[Mux.scala 27:72]
  wire  _T_2315 = _T_2281 == 4'hb; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_11; // @[el2_ifu_mem_ctl.scala 404:67]
  wire [31:0] _T_2340 = _T_2315 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2355 = _T_2354 | _T_2340; // @[Mux.scala 27:72]
  wire  _T_2318 = _T_2281 == 4'hc; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_12; // @[el2_ifu_mem_ctl.scala 403:65]
  wire [31:0] _T_2341 = _T_2318 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2356 = _T_2355 | _T_2341; // @[Mux.scala 27:72]
  wire  _T_2321 = _T_2281 == 4'hd; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_13; // @[el2_ifu_mem_ctl.scala 404:67]
  wire [31:0] _T_2342 = _T_2321 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2357 = _T_2356 | _T_2342; // @[Mux.scala 27:72]
  wire  _T_2324 = _T_2281 == 4'he; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_14; // @[el2_ifu_mem_ctl.scala 403:65]
  wire [31:0] _T_2343 = _T_2324 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2358 = _T_2357 | _T_2343; // @[Mux.scala 27:72]
  wire  _T_2327 = _T_2281 == 4'hf; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_15; // @[el2_ifu_mem_ctl.scala 404:67]
  wire [31:0] _T_2344 = _T_2327 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2359 = _T_2358 | _T_2344; // @[Mux.scala 27:72]
  wire [3:0] _T_2361 = {ifu_bus_rid_ff[2:1],_T_2240,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2362 = _T_2361 == 4'h0; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2409 = _T_2362 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2365 = _T_2361 == 4'h1; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2410 = _T_2365 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2425 = _T_2409 | _T_2410; // @[Mux.scala 27:72]
  wire  _T_2368 = _T_2361 == 4'h2; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2411 = _T_2368 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2426 = _T_2425 | _T_2411; // @[Mux.scala 27:72]
  wire  _T_2371 = _T_2361 == 4'h3; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2412 = _T_2371 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2427 = _T_2426 | _T_2412; // @[Mux.scala 27:72]
  wire  _T_2374 = _T_2361 == 4'h4; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2413 = _T_2374 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2428 = _T_2427 | _T_2413; // @[Mux.scala 27:72]
  wire  _T_2377 = _T_2361 == 4'h5; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2414 = _T_2377 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2429 = _T_2428 | _T_2414; // @[Mux.scala 27:72]
  wire  _T_2380 = _T_2361 == 4'h6; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2415 = _T_2380 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2430 = _T_2429 | _T_2415; // @[Mux.scala 27:72]
  wire  _T_2383 = _T_2361 == 4'h7; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2416 = _T_2383 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2431 = _T_2430 | _T_2416; // @[Mux.scala 27:72]
  wire  _T_2386 = _T_2361 == 4'h8; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2417 = _T_2386 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2432 = _T_2431 | _T_2417; // @[Mux.scala 27:72]
  wire  _T_2389 = _T_2361 == 4'h9; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2418 = _T_2389 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2433 = _T_2432 | _T_2418; // @[Mux.scala 27:72]
  wire  _T_2392 = _T_2361 == 4'ha; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2419 = _T_2392 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2434 = _T_2433 | _T_2419; // @[Mux.scala 27:72]
  wire  _T_2395 = _T_2361 == 4'hb; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2420 = _T_2395 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2435 = _T_2434 | _T_2420; // @[Mux.scala 27:72]
  wire  _T_2398 = _T_2361 == 4'hc; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2421 = _T_2398 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2436 = _T_2435 | _T_2421; // @[Mux.scala 27:72]
  wire  _T_2401 = _T_2361 == 4'hd; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2422 = _T_2401 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2437 = _T_2436 | _T_2422; // @[Mux.scala 27:72]
  wire  _T_2404 = _T_2361 == 4'he; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2423 = _T_2404 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2438 = _T_2437 | _T_2423; // @[Mux.scala 27:72]
  wire  _T_2407 = _T_2361 == 4'hf; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2424 = _T_2407 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2439 = _T_2438 | _T_2424; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2359,_T_2439}; // @[Cat.scala 29:58]
  wire [6:0] _T_991 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 416:13]
  wire  _T_992 = ^_T_991; // @[el2_lib.scala 416:20]
  wire [6:0] _T_998 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_1005 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 416:30]
  wire [14:0] _T_1006 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_998}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_1013 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 416:30]
  wire [30:0] _T_1022 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1013,_T_1006}; // @[el2_lib.scala 416:30]
  wire  _T_1023 = ^_T_1022; // @[el2_lib.scala 416:37]
  wire [6:0] _T_1029 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 416:47]
  wire [14:0] _T_1037 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1029}; // @[el2_lib.scala 416:47]
  wire [30:0] _T_1053 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1013,_T_1037}; // @[el2_lib.scala 416:47]
  wire  _T_1054 = ^_T_1053; // @[el2_lib.scala 416:54]
  wire [6:0] _T_1060 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 416:64]
  wire [14:0] _T_1068 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1060}; // @[el2_lib.scala 416:64]
  wire [30:0] _T_1084 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1005,_T_1068}; // @[el2_lib.scala 416:64]
  wire  _T_1085 = ^_T_1084; // @[el2_lib.scala 416:71]
  wire [7:0] _T_1092 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 416:81]
  wire [16:0] _T_1101 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1092}; // @[el2_lib.scala 416:81]
  wire [8:0] _T_1109 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 416:81]
  wire [17:0] _T_1118 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1109}; // @[el2_lib.scala 416:81]
  wire [34:0] _T_1119 = {_T_1118,_T_1101}; // @[el2_lib.scala 416:81]
  wire  _T_1120 = ^_T_1119; // @[el2_lib.scala 416:88]
  wire [7:0] _T_1127 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 416:98]
  wire [16:0] _T_1136 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1127}; // @[el2_lib.scala 416:98]
  wire [8:0] _T_1144 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 416:98]
  wire [17:0] _T_1153 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1144}; // @[el2_lib.scala 416:98]
  wire [34:0] _T_1154 = {_T_1153,_T_1136}; // @[el2_lib.scala 416:98]
  wire  _T_1155 = ^_T_1154; // @[el2_lib.scala 416:105]
  wire [7:0] _T_1162 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 416:115]
  wire [16:0] _T_1171 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_1162}; // @[el2_lib.scala 416:115]
  wire [8:0] _T_1179 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 416:115]
  wire [17:0] _T_1188 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1179}; // @[el2_lib.scala 416:115]
  wire [34:0] _T_1189 = {_T_1188,_T_1171}; // @[el2_lib.scala 416:115]
  wire  _T_1190 = ^_T_1189; // @[el2_lib.scala 416:122]
  wire [70:0] _T_1235 = {_T_570,_T_601,_T_632,_T_663,_T_698,_T_733,_T_768,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1234 = {_T_992,_T_1023,_T_1054,_T_1085,_T_1120,_T_1155,_T_1190,_T_2359,_T_2439}; // @[Cat.scala 29:58]
  wire [141:0] _T_1236 = {_T_570,_T_601,_T_632,_T_663,_T_698,_T_733,_T_768,ifu_bus_rdata_ff,_T_1234}; // @[Cat.scala 29:58]
  wire [141:0] _T_1239 = {_T_992,_T_1023,_T_1054,_T_1085,_T_1120,_T_1155,_T_1190,_T_2359,_T_2439,_T_1235}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1236 : _T_1239; // @[el2_ifu_mem_ctl.scala 360:28]
  wire  _T_1198 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 350:56]
  wire  _T_1199 = _T_1198 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 350:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 415:28]
  wire  _T_1399 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 620:35]
  wire  _T_1284 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 399:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1284; // @[el2_ifu_mem_ctl.scala 399:73]
  wire  _T_1325 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 406:118]
  wire  _T_1326 = ic_miss_buff_data_valid[0] & _T_1325; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1326; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1422 = _T_1399 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1402 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1285 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 399:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1285; // @[el2_ifu_mem_ctl.scala 399:73]
  wire  _T_1329 = ic_miss_buff_data_valid[1] & _T_1325; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1329; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1423 = _T_1402 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1430 = _T_1422 | _T_1423; // @[Mux.scala 27:72]
  wire  _T_1405 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1286 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 399:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1286; // @[el2_ifu_mem_ctl.scala 399:73]
  wire  _T_1332 = ic_miss_buff_data_valid[2] & _T_1325; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1332; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1424 = _T_1405 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1431 = _T_1430 | _T_1424; // @[Mux.scala 27:72]
  wire  _T_1408 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1287 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 399:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1287; // @[el2_ifu_mem_ctl.scala 399:73]
  wire  _T_1335 = ic_miss_buff_data_valid[3] & _T_1325; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1335; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1425 = _T_1408 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1432 = _T_1431 | _T_1425; // @[Mux.scala 27:72]
  wire  _T_1411 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1288 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 399:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 399:73]
  wire  _T_1338 = ic_miss_buff_data_valid[4] & _T_1325; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1338; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1426 = _T_1411 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1433 = _T_1432 | _T_1426; // @[Mux.scala 27:72]
  wire  _T_1414 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 399:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 399:73]
  wire  _T_1341 = ic_miss_buff_data_valid[5] & _T_1325; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1341; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1427 = _T_1414 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1434 = _T_1433 | _T_1427; // @[Mux.scala 27:72]
  wire  _T_1417 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1290 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 399:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1290; // @[el2_ifu_mem_ctl.scala 399:73]
  wire  _T_1344 = ic_miss_buff_data_valid[6] & _T_1325; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1344; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1428 = _T_1417 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1435 = _T_1434 | _T_1428; // @[Mux.scala 27:72]
  wire  _T_1420 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1291 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 399:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1291; // @[el2_ifu_mem_ctl.scala 399:73]
  wire  _T_1347 = ic_miss_buff_data_valid[7] & _T_1325; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1347; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1429 = _T_1420 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1435 | _T_1429; // @[Mux.scala 27:72]
  wire  _T_1438 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 418:58]
  wire  _T_1439 = bypass_valid_value_check & _T_1438; // @[el2_ifu_mem_ctl.scala 418:56]
  wire  _T_1441 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 418:77]
  wire  _T_1442 = _T_1439 & _T_1441; // @[el2_ifu_mem_ctl.scala 418:75]
  wire  _T_1447 = _T_1439 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 419:75]
  wire  _T_1448 = _T_1442 | _T_1447; // @[el2_ifu_mem_ctl.scala 418:95]
  wire  _T_1450 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 420:56]
  wire  _T_1453 = _T_1450 & _T_1441; // @[el2_ifu_mem_ctl.scala 420:74]
  wire  _T_1454 = _T_1448 | _T_1453; // @[el2_ifu_mem_ctl.scala 419:94]
  wire  _T_1458 = _T_1450 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 421:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 416:70]
  wire  _T_1459 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1475 = _T_1459 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1461 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1476 = _T_1461 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1483 = _T_1475 | _T_1476; // @[Mux.scala 27:72]
  wire  _T_1463 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1477 = _T_1463 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1484 = _T_1483 | _T_1477; // @[Mux.scala 27:72]
  wire  _T_1465 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1478 = _T_1465 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1485 = _T_1484 | _T_1478; // @[Mux.scala 27:72]
  wire  _T_1467 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1479 = _T_1467 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1486 = _T_1485 | _T_1479; // @[Mux.scala 27:72]
  wire  _T_1469 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1480 = _T_1469 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1487 = _T_1486 | _T_1480; // @[Mux.scala 27:72]
  wire  _T_1471 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1481 = _T_1471 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1488 = _T_1487 | _T_1481; // @[Mux.scala 27:72]
  wire  _T_1473 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1482 = _T_1473 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1489 = _T_1488 | _T_1482; // @[Mux.scala 27:72]
  wire  _T_1491 = _T_1458 & _T_1489; // @[el2_ifu_mem_ctl.scala 421:69]
  wire  _T_1492 = _T_1454 | _T_1491; // @[el2_ifu_mem_ctl.scala 420:94]
  wire [4:0] _GEN_446 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 422:95]
  wire  _T_1495 = _GEN_446 == 5'h1f; // @[el2_ifu_mem_ctl.scala 422:95]
  wire  _T_1496 = bypass_valid_value_check & _T_1495; // @[el2_ifu_mem_ctl.scala 422:56]
  wire  bypass_data_ready_in = _T_1492 | _T_1496; // @[el2_ifu_mem_ctl.scala 421:181]
  wire  _T_1497 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 426:53]
  wire  _T_1498 = _T_1497 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 426:73]
  wire  _T_1500 = _T_1498 & _T_319; // @[el2_ifu_mem_ctl.scala 426:96]
  wire  _T_1502 = _T_1500 & _T_58; // @[el2_ifu_mem_ctl.scala 426:118]
  wire  _T_1504 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 427:73]
  wire  _T_1506 = _T_1504 & _T_319; // @[el2_ifu_mem_ctl.scala 427:96]
  wire  _T_1508 = _T_1506 & _T_58; // @[el2_ifu_mem_ctl.scala 427:118]
  wire  _T_1509 = _T_1502 | _T_1508; // @[el2_ifu_mem_ctl.scala 426:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 429:58]
  wire  _T_1510 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 428:54]
  wire  _T_1511 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 428:76]
  wire  _T_1512 = _T_1510 & _T_1511; // @[el2_ifu_mem_ctl.scala 428:74]
  wire  _T_1514 = _T_1512 & _T_319; // @[el2_ifu_mem_ctl.scala 428:96]
  wire  ic_crit_wd_rdy_new_in = _T_1509 | _T_1514; // @[el2_ifu_mem_ctl.scala 427:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 630:43]
  wire  _T_1251 = ic_crit_wd_rdy | _T_2219; // @[el2_ifu_mem_ctl.scala 373:38]
  wire  _T_1253 = _T_1251 | _T_2235; // @[el2_ifu_mem_ctl.scala 373:64]
  wire  _T_1254 = ~_T_1253; // @[el2_ifu_mem_ctl.scala 373:21]
  wire  _T_1255 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 373:98]
  wire  sel_ic_data = _T_1254 & _T_1255; // @[el2_ifu_mem_ctl.scala 373:96]
  wire  _T_2442 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 473:44]
  wire  _T_1608 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 440:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 412:60]
  wire  _T_1552 = _T_1399 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1553 = _T_1402 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1560 = _T_1552 | _T_1553; // @[Mux.scala 27:72]
  wire  _T_1554 = _T_1405 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1561 = _T_1560 | _T_1554; // @[Mux.scala 27:72]
  wire  _T_1555 = _T_1408 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1562 = _T_1561 | _T_1555; // @[Mux.scala 27:72]
  wire  _T_1556 = _T_1411 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1563 = _T_1562 | _T_1556; // @[Mux.scala 27:72]
  wire  _T_1557 = _T_1414 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1564 = _T_1563 | _T_1557; // @[Mux.scala 27:72]
  wire  _T_1558 = _T_1417 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1565 = _T_1564 | _T_1558; // @[Mux.scala 27:72]
  wire  _T_1559 = _T_1420 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1565 | _T_1559; // @[Mux.scala 27:72]
  wire  _T_1591 = _T_2152 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1592 = _T_2155 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1599 = _T_1591 | _T_1592; // @[Mux.scala 27:72]
  wire  _T_1593 = _T_2158 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1600 = _T_1599 | _T_1593; // @[Mux.scala 27:72]
  wire  _T_1594 = _T_2161 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1601 = _T_1600 | _T_1594; // @[Mux.scala 27:72]
  wire  _T_1595 = _T_2164 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1602 = _T_1601 | _T_1595; // @[Mux.scala 27:72]
  wire  _T_1596 = _T_2167 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1603 = _T_1602 | _T_1596; // @[Mux.scala 27:72]
  wire  _T_1597 = _T_2170 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1604 = _T_1603 | _T_1597; // @[Mux.scala 27:72]
  wire  _T_1598 = _T_2173 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1604 | _T_1598; // @[Mux.scala 27:72]
  wire  _T_1609 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 442:70]
  wire  ifu_byp_data_err_new = _T_1608 ? ic_miss_buff_data_error_bypass : _T_1609; // @[el2_ifu_mem_ctl.scala 440:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 384:42]
  wire  _T_2443 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 473:91]
  wire  _T_2444 = ~_T_2443; // @[el2_ifu_mem_ctl.scala 473:60]
  wire  ic_rd_parity_final_err = _T_2442 & _T_2444; // @[el2_ifu_mem_ctl.scala 473:58]
  reg  ic_debug_ict_array_sel_ff; // @[el2_ifu_mem_ctl.scala 838:63]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9322 = _T_4619 & ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 765:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9324 = _T_4620 & ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9577 = _T_9322 | _T_9324; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9326 = _T_4621 & ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9578 = _T_9577 | _T_9326; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9328 = _T_4622 & ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9579 = _T_9578 | _T_9328; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9330 = _T_4623 & ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9580 = _T_9579 | _T_9330; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9332 = _T_4624 & ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9581 = _T_9580 | _T_9332; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9334 = _T_4625 & ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9582 = _T_9581 | _T_9334; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9336 = _T_4626 & ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9583 = _T_9582 | _T_9336; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9338 = _T_4627 & ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9584 = _T_9583 | _T_9338; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9340 = _T_4628 & ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9585 = _T_9584 | _T_9340; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9342 = _T_4629 & ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9586 = _T_9585 | _T_9342; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9344 = _T_4630 & ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9587 = _T_9586 | _T_9344; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9346 = _T_4631 & ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9588 = _T_9587 | _T_9346; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9348 = _T_4632 & ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9589 = _T_9588 | _T_9348; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9350 = _T_4633 & ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9590 = _T_9589 | _T_9350; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9352 = _T_4634 & ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9591 = _T_9590 | _T_9352; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9354 = _T_4635 & ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9592 = _T_9591 | _T_9354; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9356 = _T_4636 & ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9593 = _T_9592 | _T_9356; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9358 = _T_4637 & ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9594 = _T_9593 | _T_9358; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9360 = _T_4638 & ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9595 = _T_9594 | _T_9360; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9362 = _T_4639 & ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9596 = _T_9595 | _T_9362; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9364 = _T_4640 & ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9597 = _T_9596 | _T_9364; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9366 = _T_4641 & ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9598 = _T_9597 | _T_9366; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9368 = _T_4642 & ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9599 = _T_9598 | _T_9368; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9370 = _T_4643 & ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9600 = _T_9599 | _T_9370; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9372 = _T_4644 & ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9601 = _T_9600 | _T_9372; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9374 = _T_4645 & ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9602 = _T_9601 | _T_9374; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9376 = _T_4646 & ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9603 = _T_9602 | _T_9376; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9378 = _T_4647 & ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9604 = _T_9603 | _T_9378; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9380 = _T_4648 & ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9605 = _T_9604 | _T_9380; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9382 = _T_4649 & ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9606 = _T_9605 | _T_9382; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9384 = _T_4650 & ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9607 = _T_9606 | _T_9384; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9386 = _T_4651 & ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9608 = _T_9607 | _T_9386; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9388 = _T_4652 & ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9609 = _T_9608 | _T_9388; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9390 = _T_4653 & ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9610 = _T_9609 | _T_9390; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9392 = _T_4654 & ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9611 = _T_9610 | _T_9392; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9394 = _T_4655 & ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9612 = _T_9611 | _T_9394; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9396 = _T_4656 & ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9613 = _T_9612 | _T_9396; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9398 = _T_4657 & ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9614 = _T_9613 | _T_9398; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9400 = _T_4658 & ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9615 = _T_9614 | _T_9400; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9402 = _T_4659 & ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9616 = _T_9615 | _T_9402; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9404 = _T_4660 & ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9617 = _T_9616 | _T_9404; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9406 = _T_4661 & ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9618 = _T_9617 | _T_9406; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9408 = _T_4662 & ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9619 = _T_9618 | _T_9408; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9410 = _T_4663 & ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9620 = _T_9619 | _T_9410; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9412 = _T_4664 & ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9621 = _T_9620 | _T_9412; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9414 = _T_4665 & ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9622 = _T_9621 | _T_9414; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9416 = _T_4666 & ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9623 = _T_9622 | _T_9416; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9418 = _T_4667 & ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9624 = _T_9623 | _T_9418; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9420 = _T_4668 & ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9625 = _T_9624 | _T_9420; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9422 = _T_4669 & ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9626 = _T_9625 | _T_9422; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9424 = _T_4670 & ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9627 = _T_9626 | _T_9424; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9426 = _T_4671 & ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9628 = _T_9627 | _T_9426; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9428 = _T_4672 & ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9629 = _T_9628 | _T_9428; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9430 = _T_4673 & ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9630 = _T_9629 | _T_9430; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9432 = _T_4674 & ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9631 = _T_9630 | _T_9432; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9434 = _T_4675 & ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9632 = _T_9631 | _T_9434; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9436 = _T_4676 & ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9633 = _T_9632 | _T_9436; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9438 = _T_4677 & ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9634 = _T_9633 | _T_9438; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9440 = _T_4678 & ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9635 = _T_9634 | _T_9440; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9442 = _T_4679 & ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9636 = _T_9635 | _T_9442; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9444 = _T_4680 & ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9637 = _T_9636 | _T_9444; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9446 = _T_4681 & ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9638 = _T_9637 | _T_9446; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9448 = _T_4682 & ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9639 = _T_9638 | _T_9448; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9450 = _T_4683 & ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9640 = _T_9639 | _T_9450; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9452 = _T_4684 & ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9641 = _T_9640 | _T_9452; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9454 = _T_4685 & ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9642 = _T_9641 | _T_9454; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9456 = _T_4686 & ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9643 = _T_9642 | _T_9456; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9458 = _T_4687 & ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9644 = _T_9643 | _T_9458; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9460 = _T_4688 & ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9645 = _T_9644 | _T_9460; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9462 = _T_4689 & ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9646 = _T_9645 | _T_9462; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9464 = _T_4690 & ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9647 = _T_9646 | _T_9464; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9466 = _T_4691 & ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9648 = _T_9647 | _T_9466; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9468 = _T_4692 & ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9649 = _T_9648 | _T_9468; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9470 = _T_4693 & ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9650 = _T_9649 | _T_9470; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9472 = _T_4694 & ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9651 = _T_9650 | _T_9472; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9474 = _T_4695 & ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9652 = _T_9651 | _T_9474; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9476 = _T_4696 & ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9653 = _T_9652 | _T_9476; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9478 = _T_4697 & ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9654 = _T_9653 | _T_9478; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9480 = _T_4698 & ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9655 = _T_9654 | _T_9480; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9482 = _T_4699 & ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9656 = _T_9655 | _T_9482; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9484 = _T_4700 & ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9657 = _T_9656 | _T_9484; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9486 = _T_4701 & ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9658 = _T_9657 | _T_9486; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9488 = _T_4702 & ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9659 = _T_9658 | _T_9488; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9490 = _T_4703 & ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9660 = _T_9659 | _T_9490; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9492 = _T_4704 & ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9661 = _T_9660 | _T_9492; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9494 = _T_4705 & ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9662 = _T_9661 | _T_9494; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9496 = _T_4706 & ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9663 = _T_9662 | _T_9496; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9498 = _T_4707 & ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9664 = _T_9663 | _T_9498; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9500 = _T_4708 & ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9665 = _T_9664 | _T_9500; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9502 = _T_4709 & ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9666 = _T_9665 | _T_9502; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9504 = _T_4710 & ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9667 = _T_9666 | _T_9504; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9506 = _T_4711 & ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9668 = _T_9667 | _T_9506; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9508 = _T_4712 & ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9669 = _T_9668 | _T_9508; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9510 = _T_4713 & ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9670 = _T_9669 | _T_9510; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9512 = _T_4714 & ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9671 = _T_9670 | _T_9512; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9514 = _T_4715 & ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9672 = _T_9671 | _T_9514; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9516 = _T_4716 & ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9673 = _T_9672 | _T_9516; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9518 = _T_4717 & ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9674 = _T_9673 | _T_9518; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9520 = _T_4718 & ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9675 = _T_9674 | _T_9520; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9522 = _T_4719 & ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9676 = _T_9675 | _T_9522; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9524 = _T_4720 & ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9677 = _T_9676 | _T_9524; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9526 = _T_4721 & ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9678 = _T_9677 | _T_9526; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9528 = _T_4722 & ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9679 = _T_9678 | _T_9528; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9530 = _T_4723 & ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9680 = _T_9679 | _T_9530; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9532 = _T_4724 & ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9681 = _T_9680 | _T_9532; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9534 = _T_4725 & ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9682 = _T_9681 | _T_9534; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9536 = _T_4726 & ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9683 = _T_9682 | _T_9536; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9538 = _T_4727 & ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9684 = _T_9683 | _T_9538; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9540 = _T_4728 & ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9685 = _T_9684 | _T_9540; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9542 = _T_4729 & ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9686 = _T_9685 | _T_9542; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9544 = _T_4730 & ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9687 = _T_9686 | _T_9544; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9546 = _T_4731 & ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9688 = _T_9687 | _T_9546; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9548 = _T_4732 & ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9689 = _T_9688 | _T_9548; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9550 = _T_4733 & ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9690 = _T_9689 | _T_9550; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9552 = _T_4734 & ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9691 = _T_9690 | _T_9552; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9554 = _T_4735 & ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9692 = _T_9691 | _T_9554; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9556 = _T_4736 & ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9693 = _T_9692 | _T_9556; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9558 = _T_4737 & ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9694 = _T_9693 | _T_9558; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9560 = _T_4738 & ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9695 = _T_9694 | _T_9560; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9562 = _T_4739 & ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9696 = _T_9695 | _T_9562; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9564 = _T_4740 & ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9697 = _T_9696 | _T_9564; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9566 = _T_4741 & ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9698 = _T_9697 | _T_9566; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9568 = _T_4742 & ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9699 = _T_9698 | _T_9568; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9570 = _T_4743 & ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9700 = _T_9699 | _T_9570; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9572 = _T_4744 & ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9701 = _T_9700 | _T_9572; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9574 = _T_4745 & ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9702 = _T_9701 | _T_9574; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9576 = _T_4746 & ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9703 = _T_9702 | _T_9576; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_8939 = _T_4619 & ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 765:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_8941 = _T_4620 & ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9194 = _T_8939 | _T_8941; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_8943 = _T_4621 & ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9195 = _T_9194 | _T_8943; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_8945 = _T_4622 & ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9196 = _T_9195 | _T_8945; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_8947 = _T_4623 & ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9197 = _T_9196 | _T_8947; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_8949 = _T_4624 & ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9198 = _T_9197 | _T_8949; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_8951 = _T_4625 & ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9199 = _T_9198 | _T_8951; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_8953 = _T_4626 & ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9200 = _T_9199 | _T_8953; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_8955 = _T_4627 & ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9201 = _T_9200 | _T_8955; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_8957 = _T_4628 & ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9202 = _T_9201 | _T_8957; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_8959 = _T_4629 & ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9203 = _T_9202 | _T_8959; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_8961 = _T_4630 & ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9204 = _T_9203 | _T_8961; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_8963 = _T_4631 & ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9205 = _T_9204 | _T_8963; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_8965 = _T_4632 & ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9206 = _T_9205 | _T_8965; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_8967 = _T_4633 & ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9207 = _T_9206 | _T_8967; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_8969 = _T_4634 & ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9208 = _T_9207 | _T_8969; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_8971 = _T_4635 & ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9209 = _T_9208 | _T_8971; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_8973 = _T_4636 & ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9210 = _T_9209 | _T_8973; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_8975 = _T_4637 & ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9211 = _T_9210 | _T_8975; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_8977 = _T_4638 & ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9212 = _T_9211 | _T_8977; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_8979 = _T_4639 & ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9213 = _T_9212 | _T_8979; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_8981 = _T_4640 & ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9214 = _T_9213 | _T_8981; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_8983 = _T_4641 & ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9215 = _T_9214 | _T_8983; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_8985 = _T_4642 & ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9216 = _T_9215 | _T_8985; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_8987 = _T_4643 & ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9217 = _T_9216 | _T_8987; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_8989 = _T_4644 & ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9218 = _T_9217 | _T_8989; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_8991 = _T_4645 & ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9219 = _T_9218 | _T_8991; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_8993 = _T_4646 & ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9220 = _T_9219 | _T_8993; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_8995 = _T_4647 & ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9221 = _T_9220 | _T_8995; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_8997 = _T_4648 & ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9222 = _T_9221 | _T_8997; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_8999 = _T_4649 & ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9223 = _T_9222 | _T_8999; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9001 = _T_4650 & ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9224 = _T_9223 | _T_9001; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9003 = _T_4651 & ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9225 = _T_9224 | _T_9003; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9005 = _T_4652 & ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9226 = _T_9225 | _T_9005; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9007 = _T_4653 & ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9227 = _T_9226 | _T_9007; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9009 = _T_4654 & ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9228 = _T_9227 | _T_9009; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9011 = _T_4655 & ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9229 = _T_9228 | _T_9011; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9013 = _T_4656 & ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9230 = _T_9229 | _T_9013; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9015 = _T_4657 & ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9231 = _T_9230 | _T_9015; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9017 = _T_4658 & ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9232 = _T_9231 | _T_9017; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9019 = _T_4659 & ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9233 = _T_9232 | _T_9019; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9021 = _T_4660 & ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9234 = _T_9233 | _T_9021; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9023 = _T_4661 & ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9235 = _T_9234 | _T_9023; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9025 = _T_4662 & ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9236 = _T_9235 | _T_9025; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9027 = _T_4663 & ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9237 = _T_9236 | _T_9027; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9029 = _T_4664 & ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9238 = _T_9237 | _T_9029; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9031 = _T_4665 & ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9239 = _T_9238 | _T_9031; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9033 = _T_4666 & ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9240 = _T_9239 | _T_9033; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9035 = _T_4667 & ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9241 = _T_9240 | _T_9035; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9037 = _T_4668 & ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9242 = _T_9241 | _T_9037; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9039 = _T_4669 & ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9243 = _T_9242 | _T_9039; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9041 = _T_4670 & ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9244 = _T_9243 | _T_9041; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9043 = _T_4671 & ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9245 = _T_9244 | _T_9043; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9045 = _T_4672 & ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9246 = _T_9245 | _T_9045; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9047 = _T_4673 & ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9247 = _T_9246 | _T_9047; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9049 = _T_4674 & ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9248 = _T_9247 | _T_9049; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9051 = _T_4675 & ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9249 = _T_9248 | _T_9051; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9053 = _T_4676 & ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9250 = _T_9249 | _T_9053; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9055 = _T_4677 & ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9251 = _T_9250 | _T_9055; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9057 = _T_4678 & ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9252 = _T_9251 | _T_9057; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9059 = _T_4679 & ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9253 = _T_9252 | _T_9059; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9061 = _T_4680 & ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9254 = _T_9253 | _T_9061; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9063 = _T_4681 & ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9255 = _T_9254 | _T_9063; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9065 = _T_4682 & ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9256 = _T_9255 | _T_9065; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9067 = _T_4683 & ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9257 = _T_9256 | _T_9067; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9069 = _T_4684 & ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9258 = _T_9257 | _T_9069; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9071 = _T_4685 & ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9259 = _T_9258 | _T_9071; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9073 = _T_4686 & ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9260 = _T_9259 | _T_9073; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9075 = _T_4687 & ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9261 = _T_9260 | _T_9075; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9077 = _T_4688 & ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9262 = _T_9261 | _T_9077; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9079 = _T_4689 & ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9263 = _T_9262 | _T_9079; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9081 = _T_4690 & ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9264 = _T_9263 | _T_9081; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9083 = _T_4691 & ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9265 = _T_9264 | _T_9083; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9085 = _T_4692 & ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9266 = _T_9265 | _T_9085; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9087 = _T_4693 & ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9267 = _T_9266 | _T_9087; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9089 = _T_4694 & ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9268 = _T_9267 | _T_9089; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9091 = _T_4695 & ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9269 = _T_9268 | _T_9091; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9093 = _T_4696 & ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9270 = _T_9269 | _T_9093; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9095 = _T_4697 & ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9271 = _T_9270 | _T_9095; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9097 = _T_4698 & ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9272 = _T_9271 | _T_9097; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9099 = _T_4699 & ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9273 = _T_9272 | _T_9099; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9101 = _T_4700 & ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9274 = _T_9273 | _T_9101; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9103 = _T_4701 & ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9275 = _T_9274 | _T_9103; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9105 = _T_4702 & ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9276 = _T_9275 | _T_9105; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9107 = _T_4703 & ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9277 = _T_9276 | _T_9107; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9109 = _T_4704 & ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9278 = _T_9277 | _T_9109; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9111 = _T_4705 & ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9279 = _T_9278 | _T_9111; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9113 = _T_4706 & ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9280 = _T_9279 | _T_9113; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9115 = _T_4707 & ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9281 = _T_9280 | _T_9115; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9117 = _T_4708 & ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9282 = _T_9281 | _T_9117; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9119 = _T_4709 & ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9283 = _T_9282 | _T_9119; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9121 = _T_4710 & ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9284 = _T_9283 | _T_9121; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9123 = _T_4711 & ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9285 = _T_9284 | _T_9123; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9125 = _T_4712 & ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9286 = _T_9285 | _T_9125; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9127 = _T_4713 & ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9287 = _T_9286 | _T_9127; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9129 = _T_4714 & ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9288 = _T_9287 | _T_9129; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9131 = _T_4715 & ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9289 = _T_9288 | _T_9131; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9133 = _T_4716 & ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9290 = _T_9289 | _T_9133; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9135 = _T_4717 & ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9291 = _T_9290 | _T_9135; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9137 = _T_4718 & ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9292 = _T_9291 | _T_9137; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9139 = _T_4719 & ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9293 = _T_9292 | _T_9139; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9141 = _T_4720 & ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9294 = _T_9293 | _T_9141; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9143 = _T_4721 & ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9295 = _T_9294 | _T_9143; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9145 = _T_4722 & ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9296 = _T_9295 | _T_9145; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9147 = _T_4723 & ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9297 = _T_9296 | _T_9147; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9149 = _T_4724 & ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9298 = _T_9297 | _T_9149; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9151 = _T_4725 & ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9299 = _T_9298 | _T_9151; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9153 = _T_4726 & ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9300 = _T_9299 | _T_9153; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9155 = _T_4727 & ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9301 = _T_9300 | _T_9155; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9157 = _T_4728 & ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9302 = _T_9301 | _T_9157; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9159 = _T_4729 & ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9303 = _T_9302 | _T_9159; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9161 = _T_4730 & ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9304 = _T_9303 | _T_9161; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9163 = _T_4731 & ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9305 = _T_9304 | _T_9163; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9165 = _T_4732 & ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9306 = _T_9305 | _T_9165; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9167 = _T_4733 & ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9307 = _T_9306 | _T_9167; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9169 = _T_4734 & ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9308 = _T_9307 | _T_9169; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9171 = _T_4735 & ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9309 = _T_9308 | _T_9171; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9173 = _T_4736 & ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9310 = _T_9309 | _T_9173; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9175 = _T_4737 & ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9311 = _T_9310 | _T_9175; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9177 = _T_4738 & ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9312 = _T_9311 | _T_9177; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9179 = _T_4739 & ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9313 = _T_9312 | _T_9179; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9181 = _T_4740 & ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9314 = _T_9313 | _T_9181; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9183 = _T_4741 & ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9315 = _T_9314 | _T_9183; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9185 = _T_4742 & ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9316 = _T_9315 | _T_9185; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9187 = _T_4743 & ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9317 = _T_9316 | _T_9187; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9189 = _T_4744 & ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9318 = _T_9317 | _T_9189; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9191 = _T_4745 & ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9319 = _T_9318 | _T_9191; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9193 = _T_4746 & ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9320 = _T_9319 | _T_9193; // @[el2_ifu_mem_ctl.scala 765:91]
  wire [1:0] ic_tag_valid_unq = {_T_9703,_T_9320}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[el2_ifu_mem_ctl.scala 837:53]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 839:54]
  wire [1:0] _T_9743 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_9744 = ic_debug_way_ff & _T_9743; // @[el2_ifu_mem_ctl.scala 820:67]
  wire [1:0] _T_9745 = ic_tag_valid_unq & _T_9744; // @[el2_ifu_mem_ctl.scala 820:48]
  wire  ic_debug_tag_val_rd_out = |_T_9745; // @[el2_ifu_mem_ctl.scala 820:115]
  wire [70:0] _T_1210 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],6'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1211; // @[el2_ifu_mem_ctl.scala 356:63]
  wire  _T_1249 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 372:98]
  wire  sel_byp_data = _T_1253 & _T_1249; // @[el2_ifu_mem_ctl.scala 372:96]
  wire [63:0] _T_1260 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1261 = _T_1260 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 379:69]
  wire [63:0] _T_1263 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2099 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 448:31]
  wire  _T_1612 = ~ifu_fetch_addr_int_f[1]; // @[el2_ifu_mem_ctl.scala 444:38]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1613 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1661 = _T_1613 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1616 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1662 = _T_1616 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1677 = _T_1661 | _T_1662; // @[Mux.scala 27:72]
  wire  _T_1619 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1663 = _T_1619 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1678 = _T_1677 | _T_1663; // @[Mux.scala 27:72]
  wire  _T_1622 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1664 = _T_1622 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1679 = _T_1678 | _T_1664; // @[Mux.scala 27:72]
  wire  _T_1625 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1665 = _T_1625 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1680 = _T_1679 | _T_1665; // @[Mux.scala 27:72]
  wire  _T_1628 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1666 = _T_1628 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1681 = _T_1680 | _T_1666; // @[Mux.scala 27:72]
  wire  _T_1631 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1667 = _T_1631 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1682 = _T_1681 | _T_1667; // @[Mux.scala 27:72]
  wire  _T_1634 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1668 = _T_1634 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1683 = _T_1682 | _T_1668; // @[Mux.scala 27:72]
  wire  _T_1637 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1669 = _T_1637 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1684 = _T_1683 | _T_1669; // @[Mux.scala 27:72]
  wire  _T_1640 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1670 = _T_1640 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1685 = _T_1684 | _T_1670; // @[Mux.scala 27:72]
  wire  _T_1643 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1671 = _T_1643 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1686 = _T_1685 | _T_1671; // @[Mux.scala 27:72]
  wire  _T_1646 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1672 = _T_1646 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1687 = _T_1686 | _T_1672; // @[Mux.scala 27:72]
  wire  _T_1649 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1673 = _T_1649 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1688 = _T_1687 | _T_1673; // @[Mux.scala 27:72]
  wire  _T_1652 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1674 = _T_1652 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1689 = _T_1688 | _T_1674; // @[Mux.scala 27:72]
  wire  _T_1655 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1675 = _T_1655 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1690 = _T_1689 | _T_1675; // @[Mux.scala 27:72]
  wire  _T_1658 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1676 = _T_1658 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1691 = _T_1690 | _T_1676; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1693 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1741 = _T_1693 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1696 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1742 = _T_1696 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1757 = _T_1741 | _T_1742; // @[Mux.scala 27:72]
  wire  _T_1699 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1743 = _T_1699 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1758 = _T_1757 | _T_1743; // @[Mux.scala 27:72]
  wire  _T_1702 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1744 = _T_1702 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1759 = _T_1758 | _T_1744; // @[Mux.scala 27:72]
  wire  _T_1705 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1745 = _T_1705 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1760 = _T_1759 | _T_1745; // @[Mux.scala 27:72]
  wire  _T_1708 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1746 = _T_1708 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1761 = _T_1760 | _T_1746; // @[Mux.scala 27:72]
  wire  _T_1711 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1747 = _T_1711 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1762 = _T_1761 | _T_1747; // @[Mux.scala 27:72]
  wire  _T_1714 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1748 = _T_1714 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1763 = _T_1762 | _T_1748; // @[Mux.scala 27:72]
  wire  _T_1717 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1749 = _T_1717 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1764 = _T_1763 | _T_1749; // @[Mux.scala 27:72]
  wire  _T_1720 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1750 = _T_1720 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1765 = _T_1764 | _T_1750; // @[Mux.scala 27:72]
  wire  _T_1723 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1751 = _T_1723 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1766 = _T_1765 | _T_1751; // @[Mux.scala 27:72]
  wire  _T_1726 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1752 = _T_1726 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1767 = _T_1766 | _T_1752; // @[Mux.scala 27:72]
  wire  _T_1729 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1753 = _T_1729 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1768 = _T_1767 | _T_1753; // @[Mux.scala 27:72]
  wire  _T_1732 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1754 = _T_1732 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1769 = _T_1768 | _T_1754; // @[Mux.scala 27:72]
  wire  _T_1735 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1755 = _T_1735 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1770 = _T_1769 | _T_1755; // @[Mux.scala 27:72]
  wire  _T_1738 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1756 = _T_1738 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1771 = _T_1770 | _T_1756; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1773 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1821 = _T_1773 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1776 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1822 = _T_1776 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1837 = _T_1821 | _T_1822; // @[Mux.scala 27:72]
  wire  _T_1779 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1823 = _T_1779 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1838 = _T_1837 | _T_1823; // @[Mux.scala 27:72]
  wire  _T_1782 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1824 = _T_1782 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1839 = _T_1838 | _T_1824; // @[Mux.scala 27:72]
  wire  _T_1785 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1825 = _T_1785 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1840 = _T_1839 | _T_1825; // @[Mux.scala 27:72]
  wire  _T_1788 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1826 = _T_1788 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1841 = _T_1840 | _T_1826; // @[Mux.scala 27:72]
  wire  _T_1791 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1827 = _T_1791 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1842 = _T_1841 | _T_1827; // @[Mux.scala 27:72]
  wire  _T_1794 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1828 = _T_1794 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1843 = _T_1842 | _T_1828; // @[Mux.scala 27:72]
  wire  _T_1797 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1829 = _T_1797 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1844 = _T_1843 | _T_1829; // @[Mux.scala 27:72]
  wire  _T_1800 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1830 = _T_1800 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1845 = _T_1844 | _T_1830; // @[Mux.scala 27:72]
  wire  _T_1803 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1831 = _T_1803 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1846 = _T_1845 | _T_1831; // @[Mux.scala 27:72]
  wire  _T_1806 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1832 = _T_1806 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1847 = _T_1846 | _T_1832; // @[Mux.scala 27:72]
  wire  _T_1809 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1833 = _T_1809 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1848 = _T_1847 | _T_1833; // @[Mux.scala 27:72]
  wire  _T_1812 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1834 = _T_1812 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1849 = _T_1848 | _T_1834; // @[Mux.scala 27:72]
  wire  _T_1815 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1835 = _T_1815 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1850 = _T_1849 | _T_1835; // @[Mux.scala 27:72]
  wire  _T_1818 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1836 = _T_1818 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1851 = _T_1850 | _T_1836; // @[Mux.scala 27:72]
  wire [79:0] _T_1854 = {_T_1691,_T_1771,_T_1851}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1855 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1903 = _T_1855 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1858 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1904 = _T_1858 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1919 = _T_1903 | _T_1904; // @[Mux.scala 27:72]
  wire  _T_1861 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1905 = _T_1861 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1920 = _T_1919 | _T_1905; // @[Mux.scala 27:72]
  wire  _T_1864 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1906 = _T_1864 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1921 = _T_1920 | _T_1906; // @[Mux.scala 27:72]
  wire  _T_1867 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1907 = _T_1867 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1922 = _T_1921 | _T_1907; // @[Mux.scala 27:72]
  wire  _T_1870 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1908 = _T_1870 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1923 = _T_1922 | _T_1908; // @[Mux.scala 27:72]
  wire  _T_1873 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1909 = _T_1873 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1924 = _T_1923 | _T_1909; // @[Mux.scala 27:72]
  wire  _T_1876 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1910 = _T_1876 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1925 = _T_1924 | _T_1910; // @[Mux.scala 27:72]
  wire  _T_1879 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1911 = _T_1879 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1926 = _T_1925 | _T_1911; // @[Mux.scala 27:72]
  wire  _T_1882 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1912 = _T_1882 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1927 = _T_1926 | _T_1912; // @[Mux.scala 27:72]
  wire  _T_1885 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1913 = _T_1885 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1928 = _T_1927 | _T_1913; // @[Mux.scala 27:72]
  wire  _T_1888 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1914 = _T_1888 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1929 = _T_1928 | _T_1914; // @[Mux.scala 27:72]
  wire  _T_1891 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1915 = _T_1891 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1930 = _T_1929 | _T_1915; // @[Mux.scala 27:72]
  wire  _T_1894 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1916 = _T_1894 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1931 = _T_1930 | _T_1916; // @[Mux.scala 27:72]
  wire  _T_1897 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1917 = _T_1897 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1932 = _T_1931 | _T_1917; // @[Mux.scala 27:72]
  wire  _T_1900 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1918 = _T_1900 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1933 = _T_1932 | _T_1918; // @[Mux.scala 27:72]
  wire [31:0] _T_1983 = _T_1613 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1984 = _T_1616 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1983 | _T_1984; // @[Mux.scala 27:72]
  wire [31:0] _T_1985 = _T_1619 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1999 | _T_1985; // @[Mux.scala 27:72]
  wire [31:0] _T_1986 = _T_1622 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_2000 | _T_1986; // @[Mux.scala 27:72]
  wire [31:0] _T_1987 = _T_1625 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_2001 | _T_1987; // @[Mux.scala 27:72]
  wire [31:0] _T_1988 = _T_1628 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_2002 | _T_1988; // @[Mux.scala 27:72]
  wire [31:0] _T_1989 = _T_1631 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_2003 | _T_1989; // @[Mux.scala 27:72]
  wire [31:0] _T_1990 = _T_1634 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_2004 | _T_1990; // @[Mux.scala 27:72]
  wire [31:0] _T_1991 = _T_1637 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_2005 | _T_1991; // @[Mux.scala 27:72]
  wire [31:0] _T_1992 = _T_1640 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_2006 | _T_1992; // @[Mux.scala 27:72]
  wire [31:0] _T_1993 = _T_1643 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2008 = _T_2007 | _T_1993; // @[Mux.scala 27:72]
  wire [31:0] _T_1994 = _T_1646 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2009 = _T_2008 | _T_1994; // @[Mux.scala 27:72]
  wire [31:0] _T_1995 = _T_1649 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2010 = _T_2009 | _T_1995; // @[Mux.scala 27:72]
  wire [31:0] _T_1996 = _T_1652 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2011 = _T_2010 | _T_1996; // @[Mux.scala 27:72]
  wire [31:0] _T_1997 = _T_1655 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2012 = _T_2011 | _T_1997; // @[Mux.scala 27:72]
  wire [31:0] _T_1998 = _T_1658 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2013 = _T_2012 | _T_1998; // @[Mux.scala 27:72]
  wire [79:0] _T_2096 = {_T_1933,_T_2013,_T_1771}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1612 ? _T_1854 : _T_2096; // @[el2_ifu_mem_ctl.scala 444:37]
  wire [79:0] _T_2101 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2099 ? ic_byp_data_only_pre_new : _T_2101; // @[el2_ifu_mem_ctl.scala 448:30]
  wire [79:0] _GEN_447 = {{16'd0}, _T_1263}; // @[el2_ifu_mem_ctl.scala 379:114]
  wire [79:0] _T_1264 = _GEN_447 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 379:114]
  wire [79:0] _GEN_448 = {{16'd0}, _T_1261}; // @[el2_ifu_mem_ctl.scala 379:88]
  wire [79:0] ic_premux_data_temp = _GEN_448 | _T_1264; // @[el2_ifu_mem_ctl.scala 379:88]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_319; // @[el2_ifu_mem_ctl.scala 386:38]
  reg  ifc_region_acc_fault_memory_f; // @[el2_ifu_mem_ctl.scala 852:66]
  wire [1:0] _T_1272 = ifc_region_acc_fault_memory_f ? 2'h3 : 2'h0; // @[el2_ifu_mem_ctl.scala 391:10]
  wire [1:0] _T_1273 = ifc_region_acc_fault_f ? 2'h2 : _T_1272; // @[el2_ifu_mem_ctl.scala 390:8]
  wire  _T_1275 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[el2_ifu_mem_ctl.scala 392:45]
  wire  _T_1277 = byp_fetch_index == 5'h1f; // @[el2_ifu_mem_ctl.scala 392:80]
  wire  _T_1278 = ~_T_1277; // @[el2_ifu_mem_ctl.scala 392:71]
  wire  _T_1279 = _T_1275 & _T_1278; // @[el2_ifu_mem_ctl.scala 392:69]
  wire  _T_1280 = err_stop_state != 2'h2; // @[el2_ifu_mem_ctl.scala 392:131]
  wire  _T_1281 = _T_1279 & _T_1280; // @[el2_ifu_mem_ctl.scala 392:114]
  wire [6:0] _T_1353 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1}; // @[Cat.scala 29:58]
  wire  _T_1359 = ic_miss_buff_data_error[0] & _T_1325; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  _T_2640 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 626:47]
  wire  _T_2641 = _T_2640 & _T_13; // @[el2_ifu_mem_ctl.scala 626:50]
  wire  bus_ifu_wr_data_error = _T_2641 & miss_pending; // @[el2_ifu_mem_ctl.scala 626:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1359; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1363 = ic_miss_buff_data_error[1] & _T_1325; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1363; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1367 = ic_miss_buff_data_error[2] & _T_1325; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1367; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1371 = ic_miss_buff_data_error[3] & _T_1325; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1371; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1375 = ic_miss_buff_data_error[4] & _T_1325; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1375; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1379 = ic_miss_buff_data_error[5] & _T_1325; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1379; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1383 = ic_miss_buff_data_error[6] & _T_1325; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1383; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1387 = ic_miss_buff_data_error[7] & _T_1325; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1387; // @[el2_ifu_mem_ctl.scala 410:72]
  wire [6:0] _T_1393 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1}; // @[Cat.scala 29:58]
  reg [6:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2451 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2459 = _T_6 & _T_319; // @[el2_ifu_mem_ctl.scala 493:65]
  wire  _T_2460 = _T_2459 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 493:88]
  wire  _T_2462 = _T_2460 & _T_2573; // @[el2_ifu_mem_ctl.scala 493:112]
  wire  _T_2463 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2464 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 498:50]
  wire  _T_2466 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2472 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2474 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_22 = _T_2472 | _T_2474; // @[Conditional.scala 39:67]
  wire  _GEN_24 = _T_2466 ? _T_2464 : _GEN_22; // @[Conditional.scala 39:67]
  wire  _GEN_26 = _T_2463 ? _T_2464 : _GEN_24; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2451 ? _T_2462 : _GEN_26; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2451 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2465 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 499:56]
  wire  _GEN_27 = _T_2463 & _T_2465; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2451 ? 1'h0 : _GEN_27; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 484:58]
  wire  _T_2448 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 483:49]
  wire  _T_2453 = io_ic_error_start & _T_319; // @[el2_ifu_mem_ctl.scala 492:87]
  wire  _T_2467 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 502:54]
  wire  _T_2468 = _T_2467 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 502:84]
  wire  _T_2477 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 523:66]
  wire  _T_2478 = io_dec_tlu_flush_err_wb & _T_2477; // @[el2_ifu_mem_ctl.scala 523:52]
  wire  _T_2480 = _T_2478 & _T_2573; // @[el2_ifu_mem_ctl.scala 523:81]
  wire  _T_2482 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 526:59]
  wire  _T_2483 = _T_2482 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 526:86]
  wire  _T_2497 = _T_2482 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 529:81]
  wire  _T_2498 = _T_2497 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 529:103]
  wire  _T_2499 = _T_2498 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 529:126]
  wire  _T_2519 = _T_2497 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 536:103]
  wire  _T_2526 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 541:62]
  wire  _T_2527 = io_dec_tlu_flush_lower_wb & _T_2526; // @[el2_ifu_mem_ctl.scala 541:60]
  wire  _T_2528 = _T_2527 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 541:88]
  wire  _T_2529 = _T_2528 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 541:115]
  wire  _GEN_34 = _T_2525 & _T_2483; // @[Conditional.scala 39:67]
  wire  _GEN_37 = _T_2508 ? _T_2519 : _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_39 = _T_2508 | _T_2525; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_2481 ? _T_2499 : _GEN_37; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_2481 | _GEN_39; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2476 ? _T_2480 : _GEN_41; // @[Conditional.scala 40:58]
  reg  bus_cmd_req_hold; // @[el2_ifu_mem_ctl.scala 564:53]
  wire  _T_2541 = ic_act_miss_f | bus_cmd_req_hold; // @[el2_ifu_mem_ctl.scala 560:45]
  reg  ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 561:55]
  wire  _T_2542 = _T_2541 | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 560:64]
  wire  _T_2544 = _T_2542 & _T_2573; // @[el2_ifu_mem_ctl.scala 560:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2546 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 560:133]
  wire  _T_2547 = _T_2546 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 560:164]
  wire  _T_2548 = _T_2547 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 560:184]
  wire  _T_2549 = _T_2548 & miss_pending; // @[el2_ifu_mem_ctl.scala 560:204]
  wire  _T_2550 = ~_T_2549; // @[el2_ifu_mem_ctl.scala 560:112]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 592:45]
  wire  _T_2567 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 595:35]
  wire  _T_2568 = _T_2567 & miss_pending; // @[el2_ifu_mem_ctl.scala 595:53]
  wire  bus_cmd_sent = _T_2568 & _T_2573; // @[el2_ifu_mem_ctl.scala 595:68]
  wire  _T_2553 = ~bus_cmd_sent; // @[el2_ifu_mem_ctl.scala 563:61]
  wire  _T_2554 = _T_2541 & _T_2553; // @[el2_ifu_mem_ctl.scala 563:59]
  wire [2:0] _T_2558 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2560 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2562 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[el2_ifu_mem_ctl.scala 579:57]
  reg  ifu_bus_arvalid_ff; // @[el2_ifu_mem_ctl.scala 581:53]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 593:51]
  wire  _T_2588 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 603:73]
  wire  _T_2589 = _T_2574 & _T_2588; // @[el2_ifu_mem_ctl.scala 603:71]
  wire  _T_2591 = last_data_recieved_ff & _T_1325; // @[el2_ifu_mem_ctl.scala 603:114]
  wire [2:0] _T_2597 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 608:45]
  wire  _T_2601 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 611:48]
  wire  _T_2602 = _T_2601 & miss_pending; // @[el2_ifu_mem_ctl.scala 611:68]
  wire  bus_inc_cmd_beat_cnt = _T_2602 & _T_2573; // @[el2_ifu_mem_ctl.scala 611:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 613:57]
  wire  _T_2606 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 614:31]
  wire  _T_2607 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 614:71]
  wire  _T_2608 = _T_2607 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 614:87]
  wire  _T_2609 = ~_T_2608; // @[el2_ifu_mem_ctl.scala 614:55]
  wire  bus_hold_cmd_beat_cnt = _T_2606 & _T_2609; // @[el2_ifu_mem_ctl.scala 614:53]
  wire  _T_2610 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 615:46]
  wire  bus_cmd_beat_en = _T_2610 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 615:62]
  wire [2:0] _T_2613 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 617:46]
  wire [2:0] _T_2615 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2616 = bus_inc_cmd_beat_cnt ? _T_2613 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2617 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2619 = _T_2615 | _T_2616; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2619 | _T_2617; // @[Mux.scala 27:72]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 629:62]
  wire  _T_2648 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 634:50]
  wire  _T_2649 = io_ifc_dma_access_ok & _T_2648; // @[el2_ifu_mem_ctl.scala 634:47]
  wire  _T_2650 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 634:70]
  wire  _T_2654 = _T_2649 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 635:72]
  wire  _T_2655 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 635:111]
  wire  _T_2656 = _T_2654 & _T_2655; // @[el2_ifu_mem_ctl.scala 635:97]
  wire  ifc_dma_access_q_ok = _T_2656 & _T_2650; // @[el2_ifu_mem_ctl.scala 635:127]
  wire  _T_2659 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 638:40]
  wire  _T_2660 = _T_2659 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 638:58]
  wire  _T_2663 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 639:60]
  wire  _T_2664 = _T_2659 & _T_2663; // @[el2_ifu_mem_ctl.scala 639:58]
  wire  _T_2665 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 639:104]
  wire [2:0] _T_2670 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire  _T_2691 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[33]; // @[el2_lib.scala 259:74]
  wire  _T_2692 = _T_2691 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 259:74]
  wire  _T_2693 = _T_2692 ^ io_dma_mem_wdata[36]; // @[el2_lib.scala 259:74]
  wire  _T_2694 = _T_2693 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 259:74]
  wire  _T_2695 = _T_2694 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 259:74]
  wire  _T_2696 = _T_2695 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2697 = _T_2696 ^ io_dma_mem_wdata[43]; // @[el2_lib.scala 259:74]
  wire  _T_2698 = _T_2697 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 259:74]
  wire  _T_2699 = _T_2698 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 259:74]
  wire  _T_2700 = _T_2699 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2701 = _T_2700 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 259:74]
  wire  _T_2702 = _T_2701 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2703 = _T_2702 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2704 = _T_2703 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2705 = _T_2704 ^ io_dma_mem_wdata[58]; // @[el2_lib.scala 259:74]
  wire  _T_2706 = _T_2705 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 259:74]
  wire  _T_2707 = _T_2706 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 259:74]
  wire  _T_2726 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 259:74]
  wire  _T_2727 = _T_2726 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 259:74]
  wire  _T_2728 = _T_2727 ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 259:74]
  wire  _T_2729 = _T_2728 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 259:74]
  wire  _T_2730 = _T_2729 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 259:74]
  wire  _T_2731 = _T_2730 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2732 = _T_2731 ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 259:74]
  wire  _T_2733 = _T_2732 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 259:74]
  wire  _T_2734 = _T_2733 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 259:74]
  wire  _T_2735 = _T_2734 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2736 = _T_2735 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 259:74]
  wire  _T_2737 = _T_2736 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2738 = _T_2737 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2739 = _T_2738 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2740 = _T_2739 ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 259:74]
  wire  _T_2741 = _T_2740 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 259:74]
  wire  _T_2742 = _T_2741 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 259:74]
  wire  _T_2761 = io_dma_mem_wdata[33] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 259:74]
  wire  _T_2762 = _T_2761 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 259:74]
  wire  _T_2763 = _T_2762 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 259:74]
  wire  _T_2764 = _T_2763 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 259:74]
  wire  _T_2765 = _T_2764 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 259:74]
  wire  _T_2766 = _T_2765 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2767 = _T_2766 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 259:74]
  wire  _T_2768 = _T_2767 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 259:74]
  wire  _T_2769 = _T_2768 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 259:74]
  wire  _T_2770 = _T_2769 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2771 = _T_2770 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 259:74]
  wire  _T_2772 = _T_2771 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2773 = _T_2772 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2774 = _T_2773 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2775 = _T_2774 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 259:74]
  wire  _T_2776 = _T_2775 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 259:74]
  wire  _T_2777 = _T_2776 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 259:74]
  wire  _T_2793 = io_dma_mem_wdata[36] ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 259:74]
  wire  _T_2794 = _T_2793 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 259:74]
  wire  _T_2795 = _T_2794 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 259:74]
  wire  _T_2796 = _T_2795 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 259:74]
  wire  _T_2797 = _T_2796 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 259:74]
  wire  _T_2798 = _T_2797 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2799 = _T_2798 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 259:74]
  wire  _T_2800 = _T_2799 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 259:74]
  wire  _T_2801 = _T_2800 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 259:74]
  wire  _T_2802 = _T_2801 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2803 = _T_2802 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 259:74]
  wire  _T_2804 = _T_2803 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2805 = _T_2804 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2806 = _T_2805 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2822 = io_dma_mem_wdata[43] ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 259:74]
  wire  _T_2823 = _T_2822 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 259:74]
  wire  _T_2824 = _T_2823 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 259:74]
  wire  _T_2825 = _T_2824 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 259:74]
  wire  _T_2826 = _T_2825 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 259:74]
  wire  _T_2827 = _T_2826 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2828 = _T_2827 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 259:74]
  wire  _T_2829 = _T_2828 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 259:74]
  wire  _T_2830 = _T_2829 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 259:74]
  wire  _T_2831 = _T_2830 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2832 = _T_2831 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 259:74]
  wire  _T_2833 = _T_2832 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2834 = _T_2833 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2835 = _T_2834 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2842 = io_dma_mem_wdata[58] ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 259:74]
  wire  _T_2843 = _T_2842 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 259:74]
  wire  _T_2844 = _T_2843 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 259:74]
  wire  _T_2845 = _T_2844 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 259:74]
  wire  _T_2846 = _T_2845 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 259:74]
  wire [5:0] _T_2851 = {_T_2846,_T_2835,_T_2806,_T_2777,_T_2742,_T_2707}; // @[Cat.scala 29:58]
  wire  _T_2852 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 267:13]
  wire  _T_2853 = ^_T_2851; // @[el2_lib.scala 267:23]
  wire  _T_2854 = _T_2852 ^ _T_2853; // @[el2_lib.scala 267:18]
  wire  _T_2875 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[1]; // @[el2_lib.scala 259:74]
  wire  _T_2876 = _T_2875 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 259:74]
  wire  _T_2877 = _T_2876 ^ io_dma_mem_wdata[4]; // @[el2_lib.scala 259:74]
  wire  _T_2878 = _T_2877 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 259:74]
  wire  _T_2879 = _T_2878 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 259:74]
  wire  _T_2880 = _T_2879 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_2881 = _T_2880 ^ io_dma_mem_wdata[11]; // @[el2_lib.scala 259:74]
  wire  _T_2882 = _T_2881 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 259:74]
  wire  _T_2883 = _T_2882 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 259:74]
  wire  _T_2884 = _T_2883 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_2885 = _T_2884 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 259:74]
  wire  _T_2886 = _T_2885 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_2887 = _T_2886 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_2888 = _T_2887 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_2889 = _T_2888 ^ io_dma_mem_wdata[26]; // @[el2_lib.scala 259:74]
  wire  _T_2890 = _T_2889 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 259:74]
  wire  _T_2891 = _T_2890 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 259:74]
  wire  _T_2910 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 259:74]
  wire  _T_2911 = _T_2910 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 259:74]
  wire  _T_2912 = _T_2911 ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 259:74]
  wire  _T_2913 = _T_2912 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 259:74]
  wire  _T_2914 = _T_2913 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 259:74]
  wire  _T_2915 = _T_2914 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_2916 = _T_2915 ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 259:74]
  wire  _T_2917 = _T_2916 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 259:74]
  wire  _T_2918 = _T_2917 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 259:74]
  wire  _T_2919 = _T_2918 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_2920 = _T_2919 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 259:74]
  wire  _T_2921 = _T_2920 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_2922 = _T_2921 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_2923 = _T_2922 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_2924 = _T_2923 ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 259:74]
  wire  _T_2925 = _T_2924 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 259:74]
  wire  _T_2926 = _T_2925 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 259:74]
  wire  _T_2945 = io_dma_mem_wdata[1] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 259:74]
  wire  _T_2946 = _T_2945 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 259:74]
  wire  _T_2947 = _T_2946 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 259:74]
  wire  _T_2948 = _T_2947 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 259:74]
  wire  _T_2949 = _T_2948 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 259:74]
  wire  _T_2950 = _T_2949 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_2951 = _T_2950 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 259:74]
  wire  _T_2952 = _T_2951 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 259:74]
  wire  _T_2953 = _T_2952 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 259:74]
  wire  _T_2954 = _T_2953 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_2955 = _T_2954 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 259:74]
  wire  _T_2956 = _T_2955 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_2957 = _T_2956 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_2958 = _T_2957 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_2959 = _T_2958 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 259:74]
  wire  _T_2960 = _T_2959 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 259:74]
  wire  _T_2961 = _T_2960 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 259:74]
  wire  _T_2977 = io_dma_mem_wdata[4] ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 259:74]
  wire  _T_2978 = _T_2977 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 259:74]
  wire  _T_2979 = _T_2978 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 259:74]
  wire  _T_2980 = _T_2979 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 259:74]
  wire  _T_2981 = _T_2980 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 259:74]
  wire  _T_2982 = _T_2981 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_2983 = _T_2982 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 259:74]
  wire  _T_2984 = _T_2983 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 259:74]
  wire  _T_2985 = _T_2984 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 259:74]
  wire  _T_2986 = _T_2985 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_2987 = _T_2986 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 259:74]
  wire  _T_2988 = _T_2987 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_2989 = _T_2988 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_2990 = _T_2989 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_3006 = io_dma_mem_wdata[11] ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 259:74]
  wire  _T_3007 = _T_3006 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 259:74]
  wire  _T_3008 = _T_3007 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 259:74]
  wire  _T_3009 = _T_3008 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 259:74]
  wire  _T_3010 = _T_3009 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 259:74]
  wire  _T_3011 = _T_3010 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_3012 = _T_3011 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 259:74]
  wire  _T_3013 = _T_3012 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 259:74]
  wire  _T_3014 = _T_3013 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 259:74]
  wire  _T_3015 = _T_3014 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_3016 = _T_3015 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 259:74]
  wire  _T_3017 = _T_3016 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_3018 = _T_3017 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_3019 = _T_3018 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_3026 = io_dma_mem_wdata[26] ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 259:74]
  wire  _T_3027 = _T_3026 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 259:74]
  wire  _T_3028 = _T_3027 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 259:74]
  wire  _T_3029 = _T_3028 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 259:74]
  wire  _T_3030 = _T_3029 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 259:74]
  wire [5:0] _T_3035 = {_T_3030,_T_3019,_T_2990,_T_2961,_T_2926,_T_2891}; // @[Cat.scala 29:58]
  wire  _T_3036 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 267:13]
  wire  _T_3037 = ^_T_3035; // @[el2_lib.scala 267:23]
  wire  _T_3038 = _T_3036 ^ _T_3037; // @[el2_lib.scala 267:18]
  wire [6:0] _T_3039 = {_T_3038,_T_3030,_T_3019,_T_2990,_T_2961,_T_2926,_T_2891}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2854,_T_2846,_T_2835,_T_2806,_T_2777,_T_2742,_T_2707,_T_3039}; // @[Cat.scala 29:58]
  wire  _T_3041 = ~_T_2659; // @[el2_ifu_mem_ctl.scala 645:45]
  wire  _T_3042 = iccm_correct_ecc & _T_3041; // @[el2_ifu_mem_ctl.scala 645:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3043 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3050 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 659:53]
  wire  _T_3383 = _T_3295[5:0] == 6'h27; // @[el2_lib.scala 339:41]
  wire  _T_3381 = _T_3295[5:0] == 6'h26; // @[el2_lib.scala 339:41]
  wire  _T_3379 = _T_3295[5:0] == 6'h25; // @[el2_lib.scala 339:41]
  wire  _T_3377 = _T_3295[5:0] == 6'h24; // @[el2_lib.scala 339:41]
  wire  _T_3375 = _T_3295[5:0] == 6'h23; // @[el2_lib.scala 339:41]
  wire  _T_3373 = _T_3295[5:0] == 6'h22; // @[el2_lib.scala 339:41]
  wire  _T_3371 = _T_3295[5:0] == 6'h21; // @[el2_lib.scala 339:41]
  wire  _T_3369 = _T_3295[5:0] == 6'h20; // @[el2_lib.scala 339:41]
  wire  _T_3367 = _T_3295[5:0] == 6'h1f; // @[el2_lib.scala 339:41]
  wire  _T_3365 = _T_3295[5:0] == 6'h1e; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3441 = {_T_3383,_T_3381,_T_3379,_T_3377,_T_3375,_T_3373,_T_3371,_T_3369,_T_3367,_T_3365}; // @[el2_lib.scala 342:69]
  wire  _T_3363 = _T_3295[5:0] == 6'h1d; // @[el2_lib.scala 339:41]
  wire  _T_3361 = _T_3295[5:0] == 6'h1c; // @[el2_lib.scala 339:41]
  wire  _T_3359 = _T_3295[5:0] == 6'h1b; // @[el2_lib.scala 339:41]
  wire  _T_3357 = _T_3295[5:0] == 6'h1a; // @[el2_lib.scala 339:41]
  wire  _T_3355 = _T_3295[5:0] == 6'h19; // @[el2_lib.scala 339:41]
  wire  _T_3353 = _T_3295[5:0] == 6'h18; // @[el2_lib.scala 339:41]
  wire  _T_3351 = _T_3295[5:0] == 6'h17; // @[el2_lib.scala 339:41]
  wire  _T_3349 = _T_3295[5:0] == 6'h16; // @[el2_lib.scala 339:41]
  wire  _T_3347 = _T_3295[5:0] == 6'h15; // @[el2_lib.scala 339:41]
  wire  _T_3345 = _T_3295[5:0] == 6'h14; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3432 = {_T_3363,_T_3361,_T_3359,_T_3357,_T_3355,_T_3353,_T_3351,_T_3349,_T_3347,_T_3345}; // @[el2_lib.scala 342:69]
  wire  _T_3343 = _T_3295[5:0] == 6'h13; // @[el2_lib.scala 339:41]
  wire  _T_3341 = _T_3295[5:0] == 6'h12; // @[el2_lib.scala 339:41]
  wire  _T_3339 = _T_3295[5:0] == 6'h11; // @[el2_lib.scala 339:41]
  wire  _T_3337 = _T_3295[5:0] == 6'h10; // @[el2_lib.scala 339:41]
  wire  _T_3335 = _T_3295[5:0] == 6'hf; // @[el2_lib.scala 339:41]
  wire  _T_3333 = _T_3295[5:0] == 6'he; // @[el2_lib.scala 339:41]
  wire  _T_3331 = _T_3295[5:0] == 6'hd; // @[el2_lib.scala 339:41]
  wire  _T_3329 = _T_3295[5:0] == 6'hc; // @[el2_lib.scala 339:41]
  wire  _T_3327 = _T_3295[5:0] == 6'hb; // @[el2_lib.scala 339:41]
  wire  _T_3325 = _T_3295[5:0] == 6'ha; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3422 = {_T_3343,_T_3341,_T_3339,_T_3337,_T_3335,_T_3333,_T_3331,_T_3329,_T_3327,_T_3325}; // @[el2_lib.scala 342:69]
  wire  _T_3323 = _T_3295[5:0] == 6'h9; // @[el2_lib.scala 339:41]
  wire  _T_3321 = _T_3295[5:0] == 6'h8; // @[el2_lib.scala 339:41]
  wire  _T_3319 = _T_3295[5:0] == 6'h7; // @[el2_lib.scala 339:41]
  wire  _T_3317 = _T_3295[5:0] == 6'h6; // @[el2_lib.scala 339:41]
  wire  _T_3315 = _T_3295[5:0] == 6'h5; // @[el2_lib.scala 339:41]
  wire  _T_3313 = _T_3295[5:0] == 6'h4; // @[el2_lib.scala 339:41]
  wire  _T_3311 = _T_3295[5:0] == 6'h3; // @[el2_lib.scala 339:41]
  wire  _T_3309 = _T_3295[5:0] == 6'h2; // @[el2_lib.scala 339:41]
  wire  _T_3307 = _T_3295[5:0] == 6'h1; // @[el2_lib.scala 339:41]
  wire [18:0] _T_3423 = {_T_3422,_T_3323,_T_3321,_T_3319,_T_3317,_T_3315,_T_3313,_T_3311,_T_3309,_T_3307}; // @[el2_lib.scala 342:69]
  wire [38:0] _T_3443 = {_T_3441,_T_3432,_T_3423}; // @[el2_lib.scala 342:69]
  wire [7:0] _T_3398 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3404 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3398}; // @[Cat.scala 29:58]
  wire [38:0] _T_3444 = _T_3443 ^ _T_3404; // @[el2_lib.scala 342:76]
  wire [38:0] _T_3445 = _T_3299 ? _T_3444 : _T_3404; // @[el2_lib.scala 342:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3445[37:32],_T_3445[30:16],_T_3445[14:8],_T_3445[6:4],_T_3445[2]}; // @[Cat.scala 29:58]
  wire  _T_3768 = _T_3680[5:0] == 6'h27; // @[el2_lib.scala 339:41]
  wire  _T_3766 = _T_3680[5:0] == 6'h26; // @[el2_lib.scala 339:41]
  wire  _T_3764 = _T_3680[5:0] == 6'h25; // @[el2_lib.scala 339:41]
  wire  _T_3762 = _T_3680[5:0] == 6'h24; // @[el2_lib.scala 339:41]
  wire  _T_3760 = _T_3680[5:0] == 6'h23; // @[el2_lib.scala 339:41]
  wire  _T_3758 = _T_3680[5:0] == 6'h22; // @[el2_lib.scala 339:41]
  wire  _T_3756 = _T_3680[5:0] == 6'h21; // @[el2_lib.scala 339:41]
  wire  _T_3754 = _T_3680[5:0] == 6'h20; // @[el2_lib.scala 339:41]
  wire  _T_3752 = _T_3680[5:0] == 6'h1f; // @[el2_lib.scala 339:41]
  wire  _T_3750 = _T_3680[5:0] == 6'h1e; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3826 = {_T_3768,_T_3766,_T_3764,_T_3762,_T_3760,_T_3758,_T_3756,_T_3754,_T_3752,_T_3750}; // @[el2_lib.scala 342:69]
  wire  _T_3748 = _T_3680[5:0] == 6'h1d; // @[el2_lib.scala 339:41]
  wire  _T_3746 = _T_3680[5:0] == 6'h1c; // @[el2_lib.scala 339:41]
  wire  _T_3744 = _T_3680[5:0] == 6'h1b; // @[el2_lib.scala 339:41]
  wire  _T_3742 = _T_3680[5:0] == 6'h1a; // @[el2_lib.scala 339:41]
  wire  _T_3740 = _T_3680[5:0] == 6'h19; // @[el2_lib.scala 339:41]
  wire  _T_3738 = _T_3680[5:0] == 6'h18; // @[el2_lib.scala 339:41]
  wire  _T_3736 = _T_3680[5:0] == 6'h17; // @[el2_lib.scala 339:41]
  wire  _T_3734 = _T_3680[5:0] == 6'h16; // @[el2_lib.scala 339:41]
  wire  _T_3732 = _T_3680[5:0] == 6'h15; // @[el2_lib.scala 339:41]
  wire  _T_3730 = _T_3680[5:0] == 6'h14; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3817 = {_T_3748,_T_3746,_T_3744,_T_3742,_T_3740,_T_3738,_T_3736,_T_3734,_T_3732,_T_3730}; // @[el2_lib.scala 342:69]
  wire  _T_3728 = _T_3680[5:0] == 6'h13; // @[el2_lib.scala 339:41]
  wire  _T_3726 = _T_3680[5:0] == 6'h12; // @[el2_lib.scala 339:41]
  wire  _T_3724 = _T_3680[5:0] == 6'h11; // @[el2_lib.scala 339:41]
  wire  _T_3722 = _T_3680[5:0] == 6'h10; // @[el2_lib.scala 339:41]
  wire  _T_3720 = _T_3680[5:0] == 6'hf; // @[el2_lib.scala 339:41]
  wire  _T_3718 = _T_3680[5:0] == 6'he; // @[el2_lib.scala 339:41]
  wire  _T_3716 = _T_3680[5:0] == 6'hd; // @[el2_lib.scala 339:41]
  wire  _T_3714 = _T_3680[5:0] == 6'hc; // @[el2_lib.scala 339:41]
  wire  _T_3712 = _T_3680[5:0] == 6'hb; // @[el2_lib.scala 339:41]
  wire  _T_3710 = _T_3680[5:0] == 6'ha; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3807 = {_T_3728,_T_3726,_T_3724,_T_3722,_T_3720,_T_3718,_T_3716,_T_3714,_T_3712,_T_3710}; // @[el2_lib.scala 342:69]
  wire  _T_3708 = _T_3680[5:0] == 6'h9; // @[el2_lib.scala 339:41]
  wire  _T_3706 = _T_3680[5:0] == 6'h8; // @[el2_lib.scala 339:41]
  wire  _T_3704 = _T_3680[5:0] == 6'h7; // @[el2_lib.scala 339:41]
  wire  _T_3702 = _T_3680[5:0] == 6'h6; // @[el2_lib.scala 339:41]
  wire  _T_3700 = _T_3680[5:0] == 6'h5; // @[el2_lib.scala 339:41]
  wire  _T_3698 = _T_3680[5:0] == 6'h4; // @[el2_lib.scala 339:41]
  wire  _T_3696 = _T_3680[5:0] == 6'h3; // @[el2_lib.scala 339:41]
  wire  _T_3694 = _T_3680[5:0] == 6'h2; // @[el2_lib.scala 339:41]
  wire  _T_3692 = _T_3680[5:0] == 6'h1; // @[el2_lib.scala 339:41]
  wire [18:0] _T_3808 = {_T_3807,_T_3708,_T_3706,_T_3704,_T_3702,_T_3700,_T_3698,_T_3696,_T_3694,_T_3692}; // @[el2_lib.scala 342:69]
  wire [38:0] _T_3828 = {_T_3826,_T_3817,_T_3808}; // @[el2_lib.scala 342:69]
  wire [7:0] _T_3783 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3789 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3783}; // @[Cat.scala 29:58]
  wire [38:0] _T_3829 = _T_3828 ^ _T_3789; // @[el2_lib.scala 342:76]
  wire [38:0] _T_3830 = _T_3684 ? _T_3829 : _T_3789; // @[el2_lib.scala 342:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3830[37:32],_T_3830[30:16],_T_3830[14:8],_T_3830[6:4],_T_3830[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 651:35]
  wire  _T_3303 = ~_T_3295[6]; // @[el2_lib.scala 335:55]
  wire  _T_3304 = _T_3297 & _T_3303; // @[el2_lib.scala 335:53]
  wire  _T_3688 = ~_T_3680[6]; // @[el2_lib.scala 335:55]
  wire  _T_3689 = _T_3682 & _T_3688; // @[el2_lib.scala 335:53]
  wire [1:0] iccm_double_ecc_error = {_T_3304,_T_3689}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 653:53]
  wire [63:0] _T_3054 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3055 = {iccm_dma_rdata_1_muxed,_T_3445[37:32],_T_3445[30:16],_T_3445[14:8],_T_3445[6:4],_T_3445[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 655:54]
  reg [2:0] iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 656:74]
  reg  iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 661:76]
  reg  iccm_dma_ecc_error; // @[el2_ifu_mem_ctl.scala 663:74]
  reg [63:0] iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 665:75]
  wire  _T_3060 = _T_2659 & _T_2648; // @[el2_ifu_mem_ctl.scala 668:65]
  wire  _T_3064 = _T_3041 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 669:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3065 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [14:0] _T_3067 = _T_3064 ? _T_3065 : io_ifc_fetch_addr_bf[14:0]; // @[el2_ifu_mem_ctl.scala 669:8]
  wire  _T_3457 = _T_3295 == 7'h40; // @[el2_lib.scala 345:62]
  wire  _T_3458 = _T_3445[38] ^ _T_3457; // @[el2_lib.scala 345:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3458,_T_3445[31],_T_3445[15],_T_3445[7],_T_3445[3],_T_3445[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3842 = _T_3680 == 7'h40; // @[el2_lib.scala 345:62]
  wire  _T_3843 = _T_3830[38] ^ _T_3842; // @[el2_lib.scala 345:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3843,_T_3830[31],_T_3830[15],_T_3830[7],_T_3830[3],_T_3830[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3859 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 681:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 683:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 684:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 692:62]
  wire  _T_3867 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 686:76]
  wire  _T_3868 = io_iccm_rd_ecc_single_err & _T_3867; // @[el2_ifu_mem_ctl.scala 686:74]
  wire  _T_3870 = _T_3868 & _T_319; // @[el2_ifu_mem_ctl.scala 686:104]
  wire  iccm_ecc_write_status = _T_3870 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 686:127]
  wire  _T_3871 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 687:67]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 691:51]
  wire [13:0] _T_3876 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 690:102]
  wire [38:0] _T_3880 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3885 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 695:41]
  wire  _T_3886 = io_ifc_fetch_req_bf & _T_3885; // @[el2_ifu_mem_ctl.scala 695:39]
  wire  _T_3887 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 695:72]
  wire  _T_3888 = _T_3886 & _T_3887; // @[el2_ifu_mem_ctl.scala 695:70]
  wire  _T_3890 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 696:34]
  wire  _T_3891 = _T_2219 & _T_3890; // @[el2_ifu_mem_ctl.scala 696:32]
  wire  _T_3894 = _T_2235 & _T_3890; // @[el2_ifu_mem_ctl.scala 697:37]
  wire  _T_3895 = _T_3891 | _T_3894; // @[el2_ifu_mem_ctl.scala 696:88]
  wire  _T_3896 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 698:19]
  wire  _T_3898 = _T_3896 & _T_3890; // @[el2_ifu_mem_ctl.scala 698:41]
  wire  _T_3899 = _T_3895 | _T_3898; // @[el2_ifu_mem_ctl.scala 697:88]
  wire  _T_3900 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 699:19]
  wire  _T_3902 = _T_3900 & _T_3890; // @[el2_ifu_mem_ctl.scala 699:35]
  wire  _T_3903 = _T_3899 | _T_3902; // @[el2_ifu_mem_ctl.scala 698:88]
  wire  _T_3906 = _T_2234 & _T_3890; // @[el2_ifu_mem_ctl.scala 700:38]
  wire  _T_3907 = _T_3903 | _T_3906; // @[el2_ifu_mem_ctl.scala 699:88]
  wire  _T_3909 = _T_2235 & miss_state_en; // @[el2_ifu_mem_ctl.scala 701:37]
  wire  _T_3910 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 701:71]
  wire  _T_3911 = _T_3909 & _T_3910; // @[el2_ifu_mem_ctl.scala 701:54]
  wire  _T_3912 = _T_3907 | _T_3911; // @[el2_ifu_mem_ctl.scala 700:57]
  wire  _T_3913 = ~_T_3912; // @[el2_ifu_mem_ctl.scala 696:5]
  wire  _T_3914 = _T_3888 & _T_3913; // @[el2_ifu_mem_ctl.scala 695:96]
  wire  _T_3915 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 702:28]
  wire  _T_3917 = _T_3915 & _T_3885; // @[el2_ifu_mem_ctl.scala 702:50]
  wire  _T_3919 = _T_3917 & _T_3887; // @[el2_ifu_mem_ctl.scala 702:81]
  wire [1:0] _T_3922 = write_ic_16_bytes ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9728 = bus_ifu_wr_en_ff_q & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 797:74]
  wire  bus_wren_1 = _T_9728 & miss_pending; // @[el2_ifu_mem_ctl.scala 797:98]
  wire  _T_9727 = bus_ifu_wr_en_ff_q & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 797:74]
  wire  bus_wren_0 = _T_9727 & miss_pending; // @[el2_ifu_mem_ctl.scala 797:98]
  wire [1:0] bus_ic_wr_en = {bus_wren_1,bus_wren_0}; // @[Cat.scala 29:58]
  wire  _T_3928 = ~_T_108; // @[el2_ifu_mem_ctl.scala 705:106]
  wire  _T_3929 = _T_2219 & _T_3928; // @[el2_ifu_mem_ctl.scala 705:104]
  wire  _T_3930 = _T_2235 | _T_3929; // @[el2_ifu_mem_ctl.scala 705:77]
  wire  _T_3934 = ~_T_51; // @[el2_ifu_mem_ctl.scala 705:172]
  wire  _T_3935 = _T_3930 & _T_3934; // @[el2_ifu_mem_ctl.scala 705:170]
  wire  _T_3936 = ~_T_3935; // @[el2_ifu_mem_ctl.scala 705:44]
  wire  _T_3940 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 708:64]
  wire  _T_3941 = ~_T_3940; // @[el2_ifu_mem_ctl.scala 708:50]
  wire  _T_3942 = _T_276 & _T_3941; // @[el2_ifu_mem_ctl.scala 708:48]
  wire  _T_3943 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 708:81]
  wire  ic_valid = _T_3942 & _T_3943; // @[el2_ifu_mem_ctl.scala 708:79]
  wire  _T_3945 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 709:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 712:14]
  wire  _T_3948 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 715:74]
  wire  _T_9725 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 796:45]
  wire  way_status_wr_en = _T_9725 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 796:58]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 717:14]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 792:41]
  reg  way_status_new_ff; // @[el2_ifu_mem_ctl.scala 723:14]
  wire  _T_3968 = ifu_status_wr_addr_ff[2:0] == 3'h0; // @[el2_ifu_mem_ctl.scala 729:128]
  wire  _T_3969 = _T_3968 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 729:136]
  wire  _T_3972 = ifu_status_wr_addr_ff[2:0] == 3'h1; // @[el2_ifu_mem_ctl.scala 729:128]
  wire  _T_3973 = _T_3972 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 729:136]
  wire  _T_3976 = ifu_status_wr_addr_ff[2:0] == 3'h2; // @[el2_ifu_mem_ctl.scala 729:128]
  wire  _T_3977 = _T_3976 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 729:136]
  wire  _T_3980 = ifu_status_wr_addr_ff[2:0] == 3'h3; // @[el2_ifu_mem_ctl.scala 729:128]
  wire  _T_3981 = _T_3980 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 729:136]
  wire  _T_3984 = ifu_status_wr_addr_ff[2:0] == 3'h4; // @[el2_ifu_mem_ctl.scala 729:128]
  wire  _T_3985 = _T_3984 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 729:136]
  wire  _T_3988 = ifu_status_wr_addr_ff[2:0] == 3'h5; // @[el2_ifu_mem_ctl.scala 729:128]
  wire  _T_3989 = _T_3988 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 729:136]
  wire  _T_3992 = ifu_status_wr_addr_ff[2:0] == 3'h6; // @[el2_ifu_mem_ctl.scala 729:128]
  wire  _T_3993 = _T_3992 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 729:136]
  wire  _T_3996 = ifu_status_wr_addr_ff[2:0] == 3'h7; // @[el2_ifu_mem_ctl.scala 729:128]
  wire  _T_3997 = _T_3996 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 729:136]
  wire  _T_9731 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 799:84]
  wire  _T_9732 = _T_9731 & miss_pending; // @[el2_ifu_mem_ctl.scala 799:108]
  wire  bus_wren_last_1 = _T_9732 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 799:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 800:84]
  wire  _T_9734 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 801:73]
  wire  _T_9729 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 799:84]
  wire  _T_9730 = _T_9729 & miss_pending; // @[el2_ifu_mem_ctl.scala 799:108]
  wire  bus_wren_last_0 = _T_9730 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 799:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 800:84]
  wire  _T_9733 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 801:73]
  wire [1:0] ifu_tag_wren = {_T_9734,_T_9733}; // @[Cat.scala 29:58]
  wire [1:0] _T_9769 = _T_3948 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_9769 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 835:90]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 744:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 748:14]
  wire  _T_5011 = ifu_ic_rw_int_addr_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 752:78]
  wire  _T_5013 = _T_5011 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 752:87]
  wire  _T_5015 = perr_ic_index_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 753:70]
  wire  _T_5017 = _T_5015 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 753:79]
  wire  _T_5018 = _T_5013 | _T_5017; // @[el2_ifu_mem_ctl.scala 752:109]
  wire  _T_5019 = _T_5018 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 753:102]
  wire  _T_5023 = _T_5011 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 752:87]
  wire  _T_5027 = _T_5015 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 753:79]
  wire  _T_5028 = _T_5023 | _T_5027; // @[el2_ifu_mem_ctl.scala 752:109]
  wire  _T_5029 = _T_5028 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 753:102]
  wire [1:0] tag_valid_clken_0 = {_T_5029,_T_5019}; // @[Cat.scala 29:58]
  wire  _T_5031 = ifu_ic_rw_int_addr_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 752:78]
  wire  _T_5033 = _T_5031 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 752:87]
  wire  _T_5035 = perr_ic_index_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 753:70]
  wire  _T_5037 = _T_5035 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 753:79]
  wire  _T_5038 = _T_5033 | _T_5037; // @[el2_ifu_mem_ctl.scala 752:109]
  wire  _T_5039 = _T_5038 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 753:102]
  wire  _T_5043 = _T_5031 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 752:87]
  wire  _T_5047 = _T_5035 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 753:79]
  wire  _T_5048 = _T_5043 | _T_5047; // @[el2_ifu_mem_ctl.scala 752:109]
  wire  _T_5049 = _T_5048 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 753:102]
  wire [1:0] tag_valid_clken_1 = {_T_5049,_T_5039}; // @[Cat.scala 29:58]
  wire  _T_5051 = ifu_ic_rw_int_addr_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 752:78]
  wire  _T_5053 = _T_5051 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 752:87]
  wire  _T_5055 = perr_ic_index_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 753:70]
  wire  _T_5057 = _T_5055 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 753:79]
  wire  _T_5058 = _T_5053 | _T_5057; // @[el2_ifu_mem_ctl.scala 752:109]
  wire  _T_5059 = _T_5058 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 753:102]
  wire  _T_5063 = _T_5051 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 752:87]
  wire  _T_5067 = _T_5055 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 753:79]
  wire  _T_5068 = _T_5063 | _T_5067; // @[el2_ifu_mem_ctl.scala 752:109]
  wire  _T_5069 = _T_5068 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 753:102]
  wire [1:0] tag_valid_clken_2 = {_T_5069,_T_5059}; // @[Cat.scala 29:58]
  wire  _T_5071 = ifu_ic_rw_int_addr_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 752:78]
  wire  _T_5073 = _T_5071 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 752:87]
  wire  _T_5075 = perr_ic_index_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 753:70]
  wire  _T_5077 = _T_5075 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 753:79]
  wire  _T_5078 = _T_5073 | _T_5077; // @[el2_ifu_mem_ctl.scala 752:109]
  wire  _T_5079 = _T_5078 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 753:102]
  wire  _T_5083 = _T_5071 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 752:87]
  wire  _T_5087 = _T_5075 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 753:79]
  wire  _T_5088 = _T_5083 | _T_5087; // @[el2_ifu_mem_ctl.scala 752:109]
  wire  _T_5089 = _T_5088 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 753:102]
  wire [1:0] tag_valid_clken_3 = {_T_5089,_T_5079}; // @[Cat.scala 29:58]
  wire  _T_5100 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 761:97]
  wire  _T_5101 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5102 = _T_5100 & _T_5101; // @[el2_ifu_mem_ctl.scala 761:122]
  wire  _T_5105 = _T_4619 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5106 = perr_ic_index_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5108 = _T_5106 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5109 = _T_5105 | _T_5108; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5110 = _T_5109 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5120 = _T_4620 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5121 = perr_ic_index_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5123 = _T_5121 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5124 = _T_5120 | _T_5123; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5125 = _T_5124 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5135 = _T_4621 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5136 = perr_ic_index_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5138 = _T_5136 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5139 = _T_5135 | _T_5138; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5140 = _T_5139 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5150 = _T_4622 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5151 = perr_ic_index_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5153 = _T_5151 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5154 = _T_5150 | _T_5153; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5155 = _T_5154 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5165 = _T_4623 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5166 = perr_ic_index_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5168 = _T_5166 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5169 = _T_5165 | _T_5168; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5170 = _T_5169 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5180 = _T_4624 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5181 = perr_ic_index_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5183 = _T_5181 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5184 = _T_5180 | _T_5183; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5185 = _T_5184 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5195 = _T_4625 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5196 = perr_ic_index_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5198 = _T_5196 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5199 = _T_5195 | _T_5198; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5200 = _T_5199 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5210 = _T_4626 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5211 = perr_ic_index_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5213 = _T_5211 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5214 = _T_5210 | _T_5213; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5215 = _T_5214 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5225 = _T_4627 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5226 = perr_ic_index_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5228 = _T_5226 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5229 = _T_5225 | _T_5228; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5230 = _T_5229 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5240 = _T_4628 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5241 = perr_ic_index_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5243 = _T_5241 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5244 = _T_5240 | _T_5243; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5245 = _T_5244 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5255 = _T_4629 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5256 = perr_ic_index_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5258 = _T_5256 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5259 = _T_5255 | _T_5258; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5260 = _T_5259 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5270 = _T_4630 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5271 = perr_ic_index_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5273 = _T_5271 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5274 = _T_5270 | _T_5273; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5275 = _T_5274 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5285 = _T_4631 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5286 = perr_ic_index_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5288 = _T_5286 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5289 = _T_5285 | _T_5288; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5290 = _T_5289 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5300 = _T_4632 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5301 = perr_ic_index_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5303 = _T_5301 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5304 = _T_5300 | _T_5303; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5305 = _T_5304 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5315 = _T_4633 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5316 = perr_ic_index_ff == 7'he; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5318 = _T_5316 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5319 = _T_5315 | _T_5318; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5320 = _T_5319 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5330 = _T_4634 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5331 = perr_ic_index_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5333 = _T_5331 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5334 = _T_5330 | _T_5333; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5335 = _T_5334 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5345 = _T_4635 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5346 = perr_ic_index_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5348 = _T_5346 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5349 = _T_5345 | _T_5348; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5350 = _T_5349 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5360 = _T_4636 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5361 = perr_ic_index_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5363 = _T_5361 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5364 = _T_5360 | _T_5363; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5365 = _T_5364 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5375 = _T_4637 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5376 = perr_ic_index_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5378 = _T_5376 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5379 = _T_5375 | _T_5378; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5380 = _T_5379 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5390 = _T_4638 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5391 = perr_ic_index_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5393 = _T_5391 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5394 = _T_5390 | _T_5393; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5395 = _T_5394 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5405 = _T_4639 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5406 = perr_ic_index_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5408 = _T_5406 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5409 = _T_5405 | _T_5408; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5410 = _T_5409 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5420 = _T_4640 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5421 = perr_ic_index_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5423 = _T_5421 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5424 = _T_5420 | _T_5423; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5425 = _T_5424 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5435 = _T_4641 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5436 = perr_ic_index_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5438 = _T_5436 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5439 = _T_5435 | _T_5438; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5440 = _T_5439 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5450 = _T_4642 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5451 = perr_ic_index_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5453 = _T_5451 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5454 = _T_5450 | _T_5453; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5455 = _T_5454 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5465 = _T_4643 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5466 = perr_ic_index_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5468 = _T_5466 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5469 = _T_5465 | _T_5468; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5470 = _T_5469 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5480 = _T_4644 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5481 = perr_ic_index_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5483 = _T_5481 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5484 = _T_5480 | _T_5483; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5485 = _T_5484 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5495 = _T_4645 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5496 = perr_ic_index_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5498 = _T_5496 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5499 = _T_5495 | _T_5498; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5500 = _T_5499 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5510 = _T_4646 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5511 = perr_ic_index_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5513 = _T_5511 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5514 = _T_5510 | _T_5513; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5515 = _T_5514 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5525 = _T_4647 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5526 = perr_ic_index_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5528 = _T_5526 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5529 = _T_5525 | _T_5528; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5530 = _T_5529 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5540 = _T_4648 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5541 = perr_ic_index_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5543 = _T_5541 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5544 = _T_5540 | _T_5543; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5545 = _T_5544 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5555 = _T_4649 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5556 = perr_ic_index_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5558 = _T_5556 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5559 = _T_5555 | _T_5558; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5560 = _T_5559 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5570 = _T_4650 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5571 = perr_ic_index_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_5573 = _T_5571 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5574 = _T_5570 | _T_5573; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5575 = _T_5574 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5585 = _T_4619 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5588 = _T_5106 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5589 = _T_5585 | _T_5588; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5590 = _T_5589 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5600 = _T_4620 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5603 = _T_5121 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5604 = _T_5600 | _T_5603; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5605 = _T_5604 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5615 = _T_4621 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5618 = _T_5136 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5619 = _T_5615 | _T_5618; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5620 = _T_5619 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5630 = _T_4622 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5633 = _T_5151 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5634 = _T_5630 | _T_5633; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5635 = _T_5634 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5645 = _T_4623 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5648 = _T_5166 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5649 = _T_5645 | _T_5648; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5650 = _T_5649 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5660 = _T_4624 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5663 = _T_5181 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5664 = _T_5660 | _T_5663; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5665 = _T_5664 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5675 = _T_4625 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5678 = _T_5196 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5679 = _T_5675 | _T_5678; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5680 = _T_5679 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5690 = _T_4626 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5693 = _T_5211 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5694 = _T_5690 | _T_5693; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5695 = _T_5694 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5705 = _T_4627 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5708 = _T_5226 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5709 = _T_5705 | _T_5708; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5710 = _T_5709 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5720 = _T_4628 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5723 = _T_5241 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5724 = _T_5720 | _T_5723; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5725 = _T_5724 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5735 = _T_4629 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5738 = _T_5256 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5739 = _T_5735 | _T_5738; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5740 = _T_5739 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5750 = _T_4630 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5753 = _T_5271 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5754 = _T_5750 | _T_5753; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5755 = _T_5754 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5765 = _T_4631 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5768 = _T_5286 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5769 = _T_5765 | _T_5768; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5770 = _T_5769 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5780 = _T_4632 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5783 = _T_5301 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5784 = _T_5780 | _T_5783; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5785 = _T_5784 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5795 = _T_4633 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5798 = _T_5316 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5799 = _T_5795 | _T_5798; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5800 = _T_5799 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5810 = _T_4634 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5813 = _T_5331 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5814 = _T_5810 | _T_5813; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5815 = _T_5814 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5825 = _T_4635 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5828 = _T_5346 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5829 = _T_5825 | _T_5828; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5830 = _T_5829 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5840 = _T_4636 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5843 = _T_5361 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5844 = _T_5840 | _T_5843; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5845 = _T_5844 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5855 = _T_4637 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5858 = _T_5376 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5859 = _T_5855 | _T_5858; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5860 = _T_5859 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5870 = _T_4638 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5873 = _T_5391 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5874 = _T_5870 | _T_5873; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5875 = _T_5874 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5885 = _T_4639 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5888 = _T_5406 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5889 = _T_5885 | _T_5888; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5890 = _T_5889 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5900 = _T_4640 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5903 = _T_5421 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5904 = _T_5900 | _T_5903; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5905 = _T_5904 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5915 = _T_4641 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5918 = _T_5436 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5919 = _T_5915 | _T_5918; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5920 = _T_5919 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5930 = _T_4642 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5933 = _T_5451 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5934 = _T_5930 | _T_5933; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5935 = _T_5934 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5945 = _T_4643 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5948 = _T_5466 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5949 = _T_5945 | _T_5948; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5950 = _T_5949 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5960 = _T_4644 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5963 = _T_5481 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5964 = _T_5960 | _T_5963; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5965 = _T_5964 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5975 = _T_4645 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5978 = _T_5496 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5979 = _T_5975 | _T_5978; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5980 = _T_5979 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_5990 = _T_4646 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_5993 = _T_5511 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_5994 = _T_5990 | _T_5993; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_5995 = _T_5994 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6005 = _T_4647 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6008 = _T_5526 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6009 = _T_6005 | _T_6008; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6010 = _T_6009 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6020 = _T_4648 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6023 = _T_5541 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6024 = _T_6020 | _T_6023; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6025 = _T_6024 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6035 = _T_4649 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6038 = _T_5556 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6039 = _T_6035 | _T_6038; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6040 = _T_6039 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6050 = _T_4650 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6053 = _T_5571 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6054 = _T_6050 | _T_6053; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6055 = _T_6054 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6065 = _T_4651 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6066 = perr_ic_index_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6068 = _T_6066 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6069 = _T_6065 | _T_6068; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6070 = _T_6069 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6080 = _T_4652 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6081 = perr_ic_index_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6083 = _T_6081 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6084 = _T_6080 | _T_6083; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6085 = _T_6084 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6095 = _T_4653 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6096 = perr_ic_index_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6098 = _T_6096 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6099 = _T_6095 | _T_6098; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6100 = _T_6099 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6110 = _T_4654 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6111 = perr_ic_index_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6113 = _T_6111 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6114 = _T_6110 | _T_6113; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6115 = _T_6114 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6125 = _T_4655 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6126 = perr_ic_index_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6128 = _T_6126 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6129 = _T_6125 | _T_6128; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6130 = _T_6129 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6140 = _T_4656 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6141 = perr_ic_index_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6143 = _T_6141 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6144 = _T_6140 | _T_6143; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6145 = _T_6144 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6155 = _T_4657 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6156 = perr_ic_index_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6158 = _T_6156 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6159 = _T_6155 | _T_6158; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6160 = _T_6159 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6170 = _T_4658 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6171 = perr_ic_index_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6173 = _T_6171 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6174 = _T_6170 | _T_6173; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6175 = _T_6174 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6185 = _T_4659 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6186 = perr_ic_index_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6188 = _T_6186 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6189 = _T_6185 | _T_6188; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6190 = _T_6189 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6200 = _T_4660 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6201 = perr_ic_index_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6203 = _T_6201 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6204 = _T_6200 | _T_6203; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6205 = _T_6204 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6215 = _T_4661 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6216 = perr_ic_index_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6218 = _T_6216 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6219 = _T_6215 | _T_6218; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6220 = _T_6219 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6230 = _T_4662 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6231 = perr_ic_index_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6233 = _T_6231 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6234 = _T_6230 | _T_6233; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6235 = _T_6234 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6245 = _T_4663 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6246 = perr_ic_index_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6248 = _T_6246 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6249 = _T_6245 | _T_6248; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6250 = _T_6249 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6260 = _T_4664 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6261 = perr_ic_index_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6263 = _T_6261 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6264 = _T_6260 | _T_6263; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6265 = _T_6264 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6275 = _T_4665 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6276 = perr_ic_index_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6278 = _T_6276 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6279 = _T_6275 | _T_6278; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6280 = _T_6279 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6290 = _T_4666 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6291 = perr_ic_index_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6293 = _T_6291 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6294 = _T_6290 | _T_6293; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6295 = _T_6294 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6305 = _T_4667 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6306 = perr_ic_index_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6308 = _T_6306 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6309 = _T_6305 | _T_6308; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6310 = _T_6309 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6320 = _T_4668 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6321 = perr_ic_index_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6323 = _T_6321 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6324 = _T_6320 | _T_6323; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6325 = _T_6324 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6335 = _T_4669 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6336 = perr_ic_index_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6338 = _T_6336 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6339 = _T_6335 | _T_6338; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6340 = _T_6339 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6350 = _T_4670 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6351 = perr_ic_index_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6353 = _T_6351 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6354 = _T_6350 | _T_6353; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6355 = _T_6354 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6365 = _T_4671 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6366 = perr_ic_index_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6368 = _T_6366 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6369 = _T_6365 | _T_6368; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6370 = _T_6369 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6380 = _T_4672 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6381 = perr_ic_index_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6383 = _T_6381 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6384 = _T_6380 | _T_6383; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6385 = _T_6384 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6395 = _T_4673 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6396 = perr_ic_index_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6398 = _T_6396 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6399 = _T_6395 | _T_6398; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6400 = _T_6399 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6410 = _T_4674 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6411 = perr_ic_index_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6413 = _T_6411 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6414 = _T_6410 | _T_6413; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6415 = _T_6414 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6425 = _T_4675 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6426 = perr_ic_index_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6428 = _T_6426 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6429 = _T_6425 | _T_6428; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6430 = _T_6429 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6440 = _T_4676 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6441 = perr_ic_index_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6443 = _T_6441 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6444 = _T_6440 | _T_6443; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6445 = _T_6444 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6455 = _T_4677 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6456 = perr_ic_index_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6458 = _T_6456 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6459 = _T_6455 | _T_6458; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6460 = _T_6459 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6470 = _T_4678 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6471 = perr_ic_index_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6473 = _T_6471 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6474 = _T_6470 | _T_6473; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6475 = _T_6474 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6485 = _T_4679 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6486 = perr_ic_index_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6488 = _T_6486 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6489 = _T_6485 | _T_6488; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6490 = _T_6489 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6500 = _T_4680 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6501 = perr_ic_index_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6503 = _T_6501 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6504 = _T_6500 | _T_6503; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6505 = _T_6504 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6515 = _T_4681 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6516 = perr_ic_index_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6518 = _T_6516 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6519 = _T_6515 | _T_6518; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6520 = _T_6519 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6530 = _T_4682 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6531 = perr_ic_index_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_6533 = _T_6531 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6534 = _T_6530 | _T_6533; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6535 = _T_6534 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6545 = _T_4651 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6548 = _T_6066 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6549 = _T_6545 | _T_6548; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6550 = _T_6549 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6560 = _T_4652 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6563 = _T_6081 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6564 = _T_6560 | _T_6563; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6565 = _T_6564 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6575 = _T_4653 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6578 = _T_6096 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6579 = _T_6575 | _T_6578; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6580 = _T_6579 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6590 = _T_4654 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6593 = _T_6111 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6594 = _T_6590 | _T_6593; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6595 = _T_6594 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6605 = _T_4655 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6608 = _T_6126 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6609 = _T_6605 | _T_6608; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6610 = _T_6609 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6620 = _T_4656 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6623 = _T_6141 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6624 = _T_6620 | _T_6623; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6625 = _T_6624 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6635 = _T_4657 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6638 = _T_6156 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6639 = _T_6635 | _T_6638; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6640 = _T_6639 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6650 = _T_4658 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6653 = _T_6171 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6654 = _T_6650 | _T_6653; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6655 = _T_6654 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6665 = _T_4659 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6668 = _T_6186 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6669 = _T_6665 | _T_6668; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6670 = _T_6669 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6680 = _T_4660 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6683 = _T_6201 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6684 = _T_6680 | _T_6683; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6685 = _T_6684 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6695 = _T_4661 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6698 = _T_6216 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6699 = _T_6695 | _T_6698; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6700 = _T_6699 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6710 = _T_4662 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6713 = _T_6231 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6714 = _T_6710 | _T_6713; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6715 = _T_6714 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6725 = _T_4663 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6728 = _T_6246 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6729 = _T_6725 | _T_6728; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6730 = _T_6729 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6740 = _T_4664 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6743 = _T_6261 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6744 = _T_6740 | _T_6743; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6745 = _T_6744 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6755 = _T_4665 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6758 = _T_6276 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6759 = _T_6755 | _T_6758; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6760 = _T_6759 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6770 = _T_4666 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6773 = _T_6291 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6774 = _T_6770 | _T_6773; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6775 = _T_6774 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6785 = _T_4667 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6788 = _T_6306 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6789 = _T_6785 | _T_6788; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6790 = _T_6789 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6800 = _T_4668 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6803 = _T_6321 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6804 = _T_6800 | _T_6803; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6805 = _T_6804 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6815 = _T_4669 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6818 = _T_6336 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6819 = _T_6815 | _T_6818; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6820 = _T_6819 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6830 = _T_4670 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6833 = _T_6351 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6834 = _T_6830 | _T_6833; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6835 = _T_6834 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6845 = _T_4671 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6848 = _T_6366 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6849 = _T_6845 | _T_6848; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6850 = _T_6849 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6860 = _T_4672 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6863 = _T_6381 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6864 = _T_6860 | _T_6863; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6865 = _T_6864 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6875 = _T_4673 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6878 = _T_6396 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6879 = _T_6875 | _T_6878; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6880 = _T_6879 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6890 = _T_4674 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6893 = _T_6411 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6894 = _T_6890 | _T_6893; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6895 = _T_6894 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6905 = _T_4675 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6908 = _T_6426 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6909 = _T_6905 | _T_6908; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6910 = _T_6909 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6920 = _T_4676 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6923 = _T_6441 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6924 = _T_6920 | _T_6923; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6925 = _T_6924 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6935 = _T_4677 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6938 = _T_6456 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6939 = _T_6935 | _T_6938; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6940 = _T_6939 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6950 = _T_4678 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6953 = _T_6471 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6954 = _T_6950 | _T_6953; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6955 = _T_6954 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6965 = _T_4679 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6968 = _T_6486 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6969 = _T_6965 | _T_6968; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6970 = _T_6969 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6980 = _T_4680 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6983 = _T_6501 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6984 = _T_6980 | _T_6983; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_6985 = _T_6984 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_6995 = _T_4681 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_6998 = _T_6516 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_6999 = _T_6995 | _T_6998; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7000 = _T_6999 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7010 = _T_4682 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7013 = _T_6531 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7014 = _T_7010 | _T_7013; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7015 = _T_7014 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7025 = _T_4683 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7026 = perr_ic_index_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7028 = _T_7026 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7029 = _T_7025 | _T_7028; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7030 = _T_7029 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7040 = _T_4684 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7041 = perr_ic_index_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7043 = _T_7041 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7044 = _T_7040 | _T_7043; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7045 = _T_7044 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7055 = _T_4685 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7056 = perr_ic_index_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7058 = _T_7056 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7059 = _T_7055 | _T_7058; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7060 = _T_7059 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7070 = _T_4686 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7071 = perr_ic_index_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7073 = _T_7071 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7074 = _T_7070 | _T_7073; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7075 = _T_7074 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7085 = _T_4687 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7086 = perr_ic_index_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7088 = _T_7086 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7089 = _T_7085 | _T_7088; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7090 = _T_7089 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7100 = _T_4688 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7101 = perr_ic_index_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7103 = _T_7101 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7104 = _T_7100 | _T_7103; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7105 = _T_7104 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7115 = _T_4689 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7116 = perr_ic_index_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7118 = _T_7116 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7119 = _T_7115 | _T_7118; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7120 = _T_7119 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7130 = _T_4690 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7131 = perr_ic_index_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7133 = _T_7131 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7134 = _T_7130 | _T_7133; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7135 = _T_7134 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7145 = _T_4691 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7146 = perr_ic_index_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7148 = _T_7146 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7149 = _T_7145 | _T_7148; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7150 = _T_7149 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7160 = _T_4692 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7161 = perr_ic_index_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7163 = _T_7161 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7164 = _T_7160 | _T_7163; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7165 = _T_7164 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7175 = _T_4693 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7176 = perr_ic_index_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7178 = _T_7176 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7179 = _T_7175 | _T_7178; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7180 = _T_7179 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7190 = _T_4694 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7191 = perr_ic_index_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7193 = _T_7191 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7194 = _T_7190 | _T_7193; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7195 = _T_7194 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7205 = _T_4695 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7206 = perr_ic_index_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7208 = _T_7206 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7209 = _T_7205 | _T_7208; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7210 = _T_7209 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7220 = _T_4696 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7221 = perr_ic_index_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7223 = _T_7221 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7224 = _T_7220 | _T_7223; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7225 = _T_7224 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7235 = _T_4697 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7236 = perr_ic_index_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7238 = _T_7236 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7239 = _T_7235 | _T_7238; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7240 = _T_7239 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7250 = _T_4698 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7251 = perr_ic_index_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7253 = _T_7251 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7254 = _T_7250 | _T_7253; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7255 = _T_7254 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7265 = _T_4699 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7266 = perr_ic_index_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7268 = _T_7266 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7269 = _T_7265 | _T_7268; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7270 = _T_7269 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7280 = _T_4700 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7281 = perr_ic_index_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7283 = _T_7281 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7284 = _T_7280 | _T_7283; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7285 = _T_7284 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7295 = _T_4701 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7296 = perr_ic_index_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7298 = _T_7296 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7299 = _T_7295 | _T_7298; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7300 = _T_7299 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7310 = _T_4702 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7311 = perr_ic_index_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7313 = _T_7311 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7314 = _T_7310 | _T_7313; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7315 = _T_7314 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7325 = _T_4703 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7326 = perr_ic_index_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7328 = _T_7326 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7329 = _T_7325 | _T_7328; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7330 = _T_7329 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7340 = _T_4704 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7341 = perr_ic_index_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7343 = _T_7341 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7344 = _T_7340 | _T_7343; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7345 = _T_7344 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7355 = _T_4705 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7356 = perr_ic_index_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7358 = _T_7356 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7359 = _T_7355 | _T_7358; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7360 = _T_7359 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7370 = _T_4706 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7371 = perr_ic_index_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7373 = _T_7371 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7374 = _T_7370 | _T_7373; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7375 = _T_7374 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7385 = _T_4707 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7386 = perr_ic_index_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7388 = _T_7386 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7389 = _T_7385 | _T_7388; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7390 = _T_7389 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7400 = _T_4708 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7401 = perr_ic_index_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7403 = _T_7401 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7404 = _T_7400 | _T_7403; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7405 = _T_7404 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7415 = _T_4709 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7416 = perr_ic_index_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7418 = _T_7416 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7419 = _T_7415 | _T_7418; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7420 = _T_7419 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7430 = _T_4710 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7431 = perr_ic_index_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7433 = _T_7431 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7434 = _T_7430 | _T_7433; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7435 = _T_7434 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7445 = _T_4711 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7446 = perr_ic_index_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7448 = _T_7446 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7449 = _T_7445 | _T_7448; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7450 = _T_7449 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7460 = _T_4712 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7461 = perr_ic_index_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7463 = _T_7461 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7464 = _T_7460 | _T_7463; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7465 = _T_7464 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7475 = _T_4713 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7476 = perr_ic_index_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7478 = _T_7476 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7479 = _T_7475 | _T_7478; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7480 = _T_7479 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7490 = _T_4714 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7491 = perr_ic_index_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7493 = _T_7491 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7494 = _T_7490 | _T_7493; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7495 = _T_7494 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7505 = _T_4683 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7508 = _T_7026 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7509 = _T_7505 | _T_7508; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7510 = _T_7509 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7520 = _T_4684 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7523 = _T_7041 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7524 = _T_7520 | _T_7523; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7525 = _T_7524 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7535 = _T_4685 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7538 = _T_7056 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7539 = _T_7535 | _T_7538; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7540 = _T_7539 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7550 = _T_4686 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7553 = _T_7071 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7554 = _T_7550 | _T_7553; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7555 = _T_7554 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7565 = _T_4687 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7568 = _T_7086 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7569 = _T_7565 | _T_7568; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7570 = _T_7569 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7580 = _T_4688 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7583 = _T_7101 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7584 = _T_7580 | _T_7583; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7585 = _T_7584 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7595 = _T_4689 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7598 = _T_7116 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7599 = _T_7595 | _T_7598; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7600 = _T_7599 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7610 = _T_4690 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7613 = _T_7131 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7614 = _T_7610 | _T_7613; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7615 = _T_7614 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7625 = _T_4691 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7628 = _T_7146 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7629 = _T_7625 | _T_7628; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7630 = _T_7629 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7640 = _T_4692 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7643 = _T_7161 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7644 = _T_7640 | _T_7643; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7645 = _T_7644 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7655 = _T_4693 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7658 = _T_7176 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7659 = _T_7655 | _T_7658; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7660 = _T_7659 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7670 = _T_4694 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7673 = _T_7191 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7674 = _T_7670 | _T_7673; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7675 = _T_7674 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7685 = _T_4695 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7688 = _T_7206 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7689 = _T_7685 | _T_7688; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7690 = _T_7689 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7700 = _T_4696 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7703 = _T_7221 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7704 = _T_7700 | _T_7703; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7705 = _T_7704 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7715 = _T_4697 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7718 = _T_7236 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7719 = _T_7715 | _T_7718; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7720 = _T_7719 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7730 = _T_4698 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7733 = _T_7251 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7734 = _T_7730 | _T_7733; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7735 = _T_7734 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7745 = _T_4699 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7748 = _T_7266 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7749 = _T_7745 | _T_7748; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7750 = _T_7749 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7760 = _T_4700 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7763 = _T_7281 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7764 = _T_7760 | _T_7763; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7765 = _T_7764 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7775 = _T_4701 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7778 = _T_7296 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7779 = _T_7775 | _T_7778; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7780 = _T_7779 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7790 = _T_4702 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7793 = _T_7311 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7794 = _T_7790 | _T_7793; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7795 = _T_7794 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7805 = _T_4703 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7808 = _T_7326 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7809 = _T_7805 | _T_7808; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7810 = _T_7809 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7820 = _T_4704 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7823 = _T_7341 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7824 = _T_7820 | _T_7823; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7825 = _T_7824 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7835 = _T_4705 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7838 = _T_7356 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7839 = _T_7835 | _T_7838; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7840 = _T_7839 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7850 = _T_4706 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7853 = _T_7371 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7854 = _T_7850 | _T_7853; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7855 = _T_7854 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7865 = _T_4707 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7868 = _T_7386 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7869 = _T_7865 | _T_7868; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7870 = _T_7869 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7880 = _T_4708 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7883 = _T_7401 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7884 = _T_7880 | _T_7883; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7885 = _T_7884 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7895 = _T_4709 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7898 = _T_7416 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7899 = _T_7895 | _T_7898; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7900 = _T_7899 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7910 = _T_4710 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7913 = _T_7431 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7914 = _T_7910 | _T_7913; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7915 = _T_7914 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7925 = _T_4711 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7928 = _T_7446 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7929 = _T_7925 | _T_7928; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7930 = _T_7929 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7940 = _T_4712 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7943 = _T_7461 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7944 = _T_7940 | _T_7943; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7945 = _T_7944 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7955 = _T_4713 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7958 = _T_7476 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7959 = _T_7955 | _T_7958; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7960 = _T_7959 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7970 = _T_4714 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7973 = _T_7491 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7974 = _T_7970 | _T_7973; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7975 = _T_7974 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_7985 = _T_4715 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_7986 = perr_ic_index_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_7988 = _T_7986 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_7989 = _T_7985 | _T_7988; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_7990 = _T_7989 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8000 = _T_4716 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8001 = perr_ic_index_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8003 = _T_8001 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8004 = _T_8000 | _T_8003; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8005 = _T_8004 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8015 = _T_4717 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8016 = perr_ic_index_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8018 = _T_8016 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8019 = _T_8015 | _T_8018; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8020 = _T_8019 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8030 = _T_4718 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8031 = perr_ic_index_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8033 = _T_8031 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8034 = _T_8030 | _T_8033; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8035 = _T_8034 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8045 = _T_4719 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8046 = perr_ic_index_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8048 = _T_8046 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8049 = _T_8045 | _T_8048; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8050 = _T_8049 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8060 = _T_4720 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8061 = perr_ic_index_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8063 = _T_8061 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8064 = _T_8060 | _T_8063; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8065 = _T_8064 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8075 = _T_4721 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8076 = perr_ic_index_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8078 = _T_8076 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8079 = _T_8075 | _T_8078; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8080 = _T_8079 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8090 = _T_4722 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8091 = perr_ic_index_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8093 = _T_8091 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8094 = _T_8090 | _T_8093; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8095 = _T_8094 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8105 = _T_4723 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8106 = perr_ic_index_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8108 = _T_8106 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8109 = _T_8105 | _T_8108; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8110 = _T_8109 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8120 = _T_4724 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8121 = perr_ic_index_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8123 = _T_8121 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8124 = _T_8120 | _T_8123; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8125 = _T_8124 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8135 = _T_4725 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8136 = perr_ic_index_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8138 = _T_8136 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8139 = _T_8135 | _T_8138; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8140 = _T_8139 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8150 = _T_4726 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8151 = perr_ic_index_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8153 = _T_8151 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8154 = _T_8150 | _T_8153; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8155 = _T_8154 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8165 = _T_4727 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8166 = perr_ic_index_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8168 = _T_8166 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8169 = _T_8165 | _T_8168; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8170 = _T_8169 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8180 = _T_4728 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8181 = perr_ic_index_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8183 = _T_8181 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8184 = _T_8180 | _T_8183; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8185 = _T_8184 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8195 = _T_4729 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8196 = perr_ic_index_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8198 = _T_8196 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8199 = _T_8195 | _T_8198; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8200 = _T_8199 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8210 = _T_4730 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8211 = perr_ic_index_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8213 = _T_8211 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8214 = _T_8210 | _T_8213; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8215 = _T_8214 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8225 = _T_4731 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8226 = perr_ic_index_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8228 = _T_8226 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8229 = _T_8225 | _T_8228; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8230 = _T_8229 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8240 = _T_4732 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8241 = perr_ic_index_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8243 = _T_8241 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8244 = _T_8240 | _T_8243; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8245 = _T_8244 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8255 = _T_4733 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8256 = perr_ic_index_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8258 = _T_8256 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8259 = _T_8255 | _T_8258; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8260 = _T_8259 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8270 = _T_4734 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8271 = perr_ic_index_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8273 = _T_8271 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8274 = _T_8270 | _T_8273; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8275 = _T_8274 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8285 = _T_4735 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8286 = perr_ic_index_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8288 = _T_8286 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8289 = _T_8285 | _T_8288; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8290 = _T_8289 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8300 = _T_4736 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8301 = perr_ic_index_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8303 = _T_8301 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8304 = _T_8300 | _T_8303; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8305 = _T_8304 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8315 = _T_4737 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8316 = perr_ic_index_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8318 = _T_8316 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8319 = _T_8315 | _T_8318; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8320 = _T_8319 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8330 = _T_4738 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8331 = perr_ic_index_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8333 = _T_8331 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8334 = _T_8330 | _T_8333; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8335 = _T_8334 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8345 = _T_4739 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8346 = perr_ic_index_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8348 = _T_8346 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8349 = _T_8345 | _T_8348; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8350 = _T_8349 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8360 = _T_4740 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8361 = perr_ic_index_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8363 = _T_8361 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8364 = _T_8360 | _T_8363; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8365 = _T_8364 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8375 = _T_4741 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8376 = perr_ic_index_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8378 = _T_8376 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8379 = _T_8375 | _T_8378; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8380 = _T_8379 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8390 = _T_4742 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8391 = perr_ic_index_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8393 = _T_8391 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8394 = _T_8390 | _T_8393; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8395 = _T_8394 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8405 = _T_4743 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8406 = perr_ic_index_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8408 = _T_8406 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8409 = _T_8405 | _T_8408; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8410 = _T_8409 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8420 = _T_4744 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8421 = perr_ic_index_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8423 = _T_8421 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8424 = _T_8420 | _T_8423; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8425 = _T_8424 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8435 = _T_4745 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8436 = perr_ic_index_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8438 = _T_8436 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8439 = _T_8435 | _T_8438; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8440 = _T_8439 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8450 = _T_4746 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8451 = perr_ic_index_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 762:102]
  wire  _T_8453 = _T_8451 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8454 = _T_8450 | _T_8453; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8455 = _T_8454 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8465 = _T_4715 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8468 = _T_7986 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8469 = _T_8465 | _T_8468; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8470 = _T_8469 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8480 = _T_4716 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8483 = _T_8001 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8484 = _T_8480 | _T_8483; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8485 = _T_8484 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8495 = _T_4717 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8498 = _T_8016 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8499 = _T_8495 | _T_8498; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8500 = _T_8499 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8510 = _T_4718 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8513 = _T_8031 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8514 = _T_8510 | _T_8513; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8515 = _T_8514 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8525 = _T_4719 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8528 = _T_8046 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8529 = _T_8525 | _T_8528; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8530 = _T_8529 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8540 = _T_4720 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8543 = _T_8061 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8544 = _T_8540 | _T_8543; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8545 = _T_8544 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8555 = _T_4721 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8558 = _T_8076 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8559 = _T_8555 | _T_8558; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8560 = _T_8559 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8570 = _T_4722 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8573 = _T_8091 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8574 = _T_8570 | _T_8573; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8575 = _T_8574 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8585 = _T_4723 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8588 = _T_8106 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8589 = _T_8585 | _T_8588; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8590 = _T_8589 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8600 = _T_4724 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8603 = _T_8121 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8604 = _T_8600 | _T_8603; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8605 = _T_8604 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8615 = _T_4725 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8618 = _T_8136 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8619 = _T_8615 | _T_8618; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8620 = _T_8619 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8630 = _T_4726 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8633 = _T_8151 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8634 = _T_8630 | _T_8633; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8635 = _T_8634 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8645 = _T_4727 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8648 = _T_8166 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8649 = _T_8645 | _T_8648; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8650 = _T_8649 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8660 = _T_4728 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8663 = _T_8181 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8664 = _T_8660 | _T_8663; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8665 = _T_8664 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8675 = _T_4729 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8678 = _T_8196 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8679 = _T_8675 | _T_8678; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8680 = _T_8679 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8690 = _T_4730 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8693 = _T_8211 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8694 = _T_8690 | _T_8693; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8695 = _T_8694 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8705 = _T_4731 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8708 = _T_8226 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8709 = _T_8705 | _T_8708; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8710 = _T_8709 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8720 = _T_4732 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8723 = _T_8241 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8724 = _T_8720 | _T_8723; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8725 = _T_8724 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8735 = _T_4733 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8738 = _T_8256 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8739 = _T_8735 | _T_8738; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8740 = _T_8739 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8750 = _T_4734 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8753 = _T_8271 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8754 = _T_8750 | _T_8753; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8755 = _T_8754 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8765 = _T_4735 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8768 = _T_8286 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8769 = _T_8765 | _T_8768; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8770 = _T_8769 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8780 = _T_4736 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8783 = _T_8301 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8784 = _T_8780 | _T_8783; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8785 = _T_8784 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8795 = _T_4737 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8798 = _T_8316 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8799 = _T_8795 | _T_8798; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8800 = _T_8799 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8810 = _T_4738 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8813 = _T_8331 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8814 = _T_8810 | _T_8813; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8815 = _T_8814 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8825 = _T_4739 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8828 = _T_8346 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8829 = _T_8825 | _T_8828; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8830 = _T_8829 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8840 = _T_4740 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8843 = _T_8361 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8844 = _T_8840 | _T_8843; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8845 = _T_8844 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8855 = _T_4741 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8858 = _T_8376 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8859 = _T_8855 | _T_8858; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8860 = _T_8859 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8870 = _T_4742 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8873 = _T_8391 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8874 = _T_8870 | _T_8873; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8875 = _T_8874 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8885 = _T_4743 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8888 = _T_8406 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8889 = _T_8885 | _T_8888; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8890 = _T_8889 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8900 = _T_4744 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8903 = _T_8421 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8904 = _T_8900 | _T_8903; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8905 = _T_8904 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8915 = _T_4745 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8918 = _T_8436 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8919 = _T_8915 | _T_8918; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8920 = _T_8919 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_8930 = _T_4746 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:59]
  wire  _T_8933 = _T_8451 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 762:124]
  wire  _T_8934 = _T_8930 | _T_8933; // @[el2_ifu_mem_ctl.scala 762:81]
  wire  _T_8935 = _T_8934 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 762:147]
  wire  _T_9737 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 817:63]
  wire  _T_9738 = _T_9737 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 817:85]
  wire [1:0] _T_9740 = _T_9738 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_9747; // @[el2_ifu_mem_ctl.scala 822:57]
  reg  _T_9748; // @[el2_ifu_mem_ctl.scala 823:56]
  reg  _T_9749; // @[el2_ifu_mem_ctl.scala 824:59]
  wire  _T_9750 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 825:80]
  wire  _T_9751 = ifu_bus_arvalid_ff & _T_9750; // @[el2_ifu_mem_ctl.scala 825:78]
  reg  _T_9753; // @[el2_ifu_mem_ctl.scala 825:58]
  reg  _T_9754; // @[el2_ifu_mem_ctl.scala 826:58]
  wire  _T_9757 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 833:71]
  wire  _T_9759 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 833:124]
  wire  _T_9761 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 834:50]
  wire  _T_9763 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 834:103]
  wire [3:0] _T_9766 = {_T_9757,_T_9759,_T_9761,_T_9763}; // @[Cat.scala 29:58]
  reg  _T_9775; // @[Reg.scala 27:20]
  wire [31:0] _T_9785 = {io_ifc_fetch_addr_bf,1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_9786 = _T_9785 | 32'h7fffffff; // @[el2_ifu_mem_ctl.scala 842:65]
  wire  _T_9788 = _T_9786 == 32'h7fffffff; // @[el2_ifu_mem_ctl.scala 842:96]
  wire [31:0] _T_9792 = _T_9785 | 32'h3fffffff; // @[el2_ifu_mem_ctl.scala 843:65]
  wire  _T_9794 = _T_9792 == 32'hffffffff; // @[el2_ifu_mem_ctl.scala 843:96]
  wire  _T_9796 = _T_9788 | _T_9794; // @[el2_ifu_mem_ctl.scala 842:162]
  wire [31:0] _T_9798 = _T_9785 | 32'h1fffffff; // @[el2_ifu_mem_ctl.scala 844:65]
  wire  _T_9800 = _T_9798 == 32'hbfffffff; // @[el2_ifu_mem_ctl.scala 844:96]
  wire  _T_9802 = _T_9796 | _T_9800; // @[el2_ifu_mem_ctl.scala 843:162]
  wire [31:0] _T_9804 = _T_9785 | 32'hfffffff; // @[el2_ifu_mem_ctl.scala 845:65]
  wire  _T_9806 = _T_9804 == 32'h8fffffff; // @[el2_ifu_mem_ctl.scala 845:96]
  wire  ifc_region_acc_okay = _T_9802 | _T_9806; // @[el2_ifu_mem_ctl.scala 844:162]
  wire  _T_9833 = ~ifc_region_acc_okay; // @[el2_ifu_mem_ctl.scala 850:65]
  wire  _T_9834 = _T_3887 & _T_9833; // @[el2_ifu_mem_ctl.scala 850:63]
  wire  ifc_region_acc_fault_memory_bf = _T_9834 & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 850:86]
  rvclkhdr rvclkhdr ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  rvclkhdr rvclkhdr_26 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_26_io_l1clk),
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en),
    .io_scan_mode(rvclkhdr_26_io_scan_mode)
  );
  rvclkhdr rvclkhdr_27 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_27_io_l1clk),
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en),
    .io_scan_mode(rvclkhdr_27_io_scan_mode)
  );
  rvclkhdr rvclkhdr_28 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_28_io_l1clk),
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en),
    .io_scan_mode(rvclkhdr_28_io_scan_mode)
  );
  rvclkhdr rvclkhdr_29 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_29_io_l1clk),
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en),
    .io_scan_mode(rvclkhdr_29_io_scan_mode)
  );
  rvclkhdr rvclkhdr_30 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_30_io_l1clk),
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en),
    .io_scan_mode(rvclkhdr_30_io_scan_mode)
  );
  rvclkhdr rvclkhdr_31 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_31_io_l1clk),
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en),
    .io_scan_mode(rvclkhdr_31_io_scan_mode)
  );
  rvclkhdr rvclkhdr_32 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_32_io_l1clk),
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en),
    .io_scan_mode(rvclkhdr_32_io_scan_mode)
  );
  rvclkhdr rvclkhdr_33 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_33_io_l1clk),
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en),
    .io_scan_mode(rvclkhdr_33_io_scan_mode)
  );
  rvclkhdr rvclkhdr_34 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_34_io_l1clk),
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en),
    .io_scan_mode(rvclkhdr_34_io_scan_mode)
  );
  rvclkhdr rvclkhdr_35 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_35_io_l1clk),
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en),
    .io_scan_mode(rvclkhdr_35_io_scan_mode)
  );
  rvclkhdr rvclkhdr_36 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_36_io_l1clk),
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en),
    .io_scan_mode(rvclkhdr_36_io_scan_mode)
  );
  rvclkhdr rvclkhdr_37 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_37_io_l1clk),
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en),
    .io_scan_mode(rvclkhdr_37_io_scan_mode)
  );
  rvclkhdr rvclkhdr_38 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_38_io_l1clk),
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en),
    .io_scan_mode(rvclkhdr_38_io_scan_mode)
  );
  rvclkhdr rvclkhdr_39 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_39_io_l1clk),
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en),
    .io_scan_mode(rvclkhdr_39_io_scan_mode)
  );
  rvclkhdr rvclkhdr_40 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_40_io_l1clk),
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en),
    .io_scan_mode(rvclkhdr_40_io_scan_mode)
  );
  rvclkhdr rvclkhdr_41 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_41_io_l1clk),
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en),
    .io_scan_mode(rvclkhdr_41_io_scan_mode)
  );
  rvclkhdr rvclkhdr_42 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_42_io_l1clk),
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en),
    .io_scan_mode(rvclkhdr_42_io_scan_mode)
  );
  rvclkhdr rvclkhdr_43 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_43_io_l1clk),
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en),
    .io_scan_mode(rvclkhdr_43_io_scan_mode)
  );
  rvclkhdr rvclkhdr_44 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_44_io_l1clk),
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en),
    .io_scan_mode(rvclkhdr_44_io_scan_mode)
  );
  rvclkhdr rvclkhdr_45 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_45_io_l1clk),
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en),
    .io_scan_mode(rvclkhdr_45_io_scan_mode)
  );
  rvclkhdr rvclkhdr_46 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_46_io_l1clk),
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en),
    .io_scan_mode(rvclkhdr_46_io_scan_mode)
  );
  rvclkhdr rvclkhdr_47 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_47_io_l1clk),
    .io_clk(rvclkhdr_47_io_clk),
    .io_en(rvclkhdr_47_io_en),
    .io_scan_mode(rvclkhdr_47_io_scan_mode)
  );
  rvclkhdr rvclkhdr_48 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_48_io_l1clk),
    .io_clk(rvclkhdr_48_io_clk),
    .io_en(rvclkhdr_48_io_en),
    .io_scan_mode(rvclkhdr_48_io_scan_mode)
  );
  rvclkhdr rvclkhdr_49 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_49_io_l1clk),
    .io_clk(rvclkhdr_49_io_clk),
    .io_en(rvclkhdr_49_io_en),
    .io_scan_mode(rvclkhdr_49_io_scan_mode)
  );
  rvclkhdr rvclkhdr_50 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_50_io_l1clk),
    .io_clk(rvclkhdr_50_io_clk),
    .io_en(rvclkhdr_50_io_en),
    .io_scan_mode(rvclkhdr_50_io_scan_mode)
  );
  rvclkhdr rvclkhdr_51 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_51_io_l1clk),
    .io_clk(rvclkhdr_51_io_clk),
    .io_en(rvclkhdr_51_io_en),
    .io_scan_mode(rvclkhdr_51_io_scan_mode)
  );
  rvclkhdr rvclkhdr_52 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_52_io_l1clk),
    .io_clk(rvclkhdr_52_io_clk),
    .io_en(rvclkhdr_52_io_en),
    .io_scan_mode(rvclkhdr_52_io_scan_mode)
  );
  rvclkhdr rvclkhdr_53 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_53_io_l1clk),
    .io_clk(rvclkhdr_53_io_clk),
    .io_en(rvclkhdr_53_io_en),
    .io_scan_mode(rvclkhdr_53_io_scan_mode)
  );
  rvclkhdr rvclkhdr_54 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_54_io_l1clk),
    .io_clk(rvclkhdr_54_io_clk),
    .io_en(rvclkhdr_54_io_en),
    .io_scan_mode(rvclkhdr_54_io_scan_mode)
  );
  rvclkhdr rvclkhdr_55 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_55_io_l1clk),
    .io_clk(rvclkhdr_55_io_clk),
    .io_en(rvclkhdr_55_io_en),
    .io_scan_mode(rvclkhdr_55_io_scan_mode)
  );
  rvclkhdr rvclkhdr_56 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_56_io_l1clk),
    .io_clk(rvclkhdr_56_io_clk),
    .io_en(rvclkhdr_56_io_en),
    .io_scan_mode(rvclkhdr_56_io_scan_mode)
  );
  rvclkhdr rvclkhdr_57 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_57_io_l1clk),
    .io_clk(rvclkhdr_57_io_clk),
    .io_en(rvclkhdr_57_io_en),
    .io_scan_mode(rvclkhdr_57_io_scan_mode)
  );
  rvclkhdr rvclkhdr_58 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_58_io_l1clk),
    .io_clk(rvclkhdr_58_io_clk),
    .io_en(rvclkhdr_58_io_en),
    .io_scan_mode(rvclkhdr_58_io_scan_mode)
  );
  rvclkhdr rvclkhdr_59 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_59_io_l1clk),
    .io_clk(rvclkhdr_59_io_clk),
    .io_en(rvclkhdr_59_io_en),
    .io_scan_mode(rvclkhdr_59_io_scan_mode)
  );
  rvclkhdr rvclkhdr_60 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_60_io_l1clk),
    .io_clk(rvclkhdr_60_io_clk),
    .io_en(rvclkhdr_60_io_en),
    .io_scan_mode(rvclkhdr_60_io_scan_mode)
  );
  rvclkhdr rvclkhdr_61 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_61_io_l1clk),
    .io_clk(rvclkhdr_61_io_clk),
    .io_en(rvclkhdr_61_io_en),
    .io_scan_mode(rvclkhdr_61_io_scan_mode)
  );
  rvclkhdr rvclkhdr_62 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_62_io_l1clk),
    .io_clk(rvclkhdr_62_io_clk),
    .io_en(rvclkhdr_62_io_en),
    .io_scan_mode(rvclkhdr_62_io_scan_mode)
  );
  rvclkhdr rvclkhdr_63 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_63_io_l1clk),
    .io_clk(rvclkhdr_63_io_clk),
    .io_en(rvclkhdr_63_io_en),
    .io_scan_mode(rvclkhdr_63_io_scan_mode)
  );
  rvclkhdr rvclkhdr_64 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_64_io_l1clk),
    .io_clk(rvclkhdr_64_io_clk),
    .io_en(rvclkhdr_64_io_en),
    .io_scan_mode(rvclkhdr_64_io_scan_mode)
  );
  rvclkhdr rvclkhdr_65 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_65_io_l1clk),
    .io_clk(rvclkhdr_65_io_clk),
    .io_en(rvclkhdr_65_io_en),
    .io_scan_mode(rvclkhdr_65_io_scan_mode)
  );
  rvclkhdr rvclkhdr_66 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_66_io_l1clk),
    .io_clk(rvclkhdr_66_io_clk),
    .io_en(rvclkhdr_66_io_en),
    .io_scan_mode(rvclkhdr_66_io_scan_mode)
  );
  rvclkhdr rvclkhdr_67 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_67_io_l1clk),
    .io_clk(rvclkhdr_67_io_clk),
    .io_en(rvclkhdr_67_io_en),
    .io_scan_mode(rvclkhdr_67_io_scan_mode)
  );
  rvclkhdr rvclkhdr_68 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_68_io_l1clk),
    .io_clk(rvclkhdr_68_io_clk),
    .io_en(rvclkhdr_68_io_en),
    .io_scan_mode(rvclkhdr_68_io_scan_mode)
  );
  rvclkhdr rvclkhdr_69 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_69_io_l1clk),
    .io_clk(rvclkhdr_69_io_clk),
    .io_en(rvclkhdr_69_io_en),
    .io_scan_mode(rvclkhdr_69_io_scan_mode)
  );
  rvclkhdr rvclkhdr_70 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_70_io_l1clk),
    .io_clk(rvclkhdr_70_io_clk),
    .io_en(rvclkhdr_70_io_en),
    .io_scan_mode(rvclkhdr_70_io_scan_mode)
  );
  rvclkhdr rvclkhdr_71 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_71_io_l1clk),
    .io_clk(rvclkhdr_71_io_clk),
    .io_en(rvclkhdr_71_io_en),
    .io_scan_mode(rvclkhdr_71_io_scan_mode)
  );
  rvclkhdr rvclkhdr_72 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_72_io_l1clk),
    .io_clk(rvclkhdr_72_io_clk),
    .io_en(rvclkhdr_72_io_en),
    .io_scan_mode(rvclkhdr_72_io_scan_mode)
  );
  rvclkhdr rvclkhdr_73 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_73_io_l1clk),
    .io_clk(rvclkhdr_73_io_clk),
    .io_en(rvclkhdr_73_io_en),
    .io_scan_mode(rvclkhdr_73_io_scan_mode)
  );
  rvclkhdr rvclkhdr_74 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_74_io_l1clk),
    .io_clk(rvclkhdr_74_io_clk),
    .io_en(rvclkhdr_74_io_en),
    .io_scan_mode(rvclkhdr_74_io_scan_mode)
  );
  rvclkhdr rvclkhdr_75 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_75_io_l1clk),
    .io_clk(rvclkhdr_75_io_clk),
    .io_en(rvclkhdr_75_io_en),
    .io_scan_mode(rvclkhdr_75_io_scan_mode)
  );
  rvclkhdr rvclkhdr_76 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_76_io_l1clk),
    .io_clk(rvclkhdr_76_io_clk),
    .io_en(rvclkhdr_76_io_en),
    .io_scan_mode(rvclkhdr_76_io_scan_mode)
  );
  rvclkhdr rvclkhdr_77 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_77_io_l1clk),
    .io_clk(rvclkhdr_77_io_clk),
    .io_en(rvclkhdr_77_io_en),
    .io_scan_mode(rvclkhdr_77_io_scan_mode)
  );
  rvclkhdr rvclkhdr_78 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_78_io_l1clk),
    .io_clk(rvclkhdr_78_io_clk),
    .io_en(rvclkhdr_78_io_en),
    .io_scan_mode(rvclkhdr_78_io_scan_mode)
  );
  rvclkhdr rvclkhdr_79 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_79_io_l1clk),
    .io_clk(rvclkhdr_79_io_clk),
    .io_en(rvclkhdr_79_io_en),
    .io_scan_mode(rvclkhdr_79_io_scan_mode)
  );
  rvclkhdr rvclkhdr_80 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_80_io_l1clk),
    .io_clk(rvclkhdr_80_io_clk),
    .io_en(rvclkhdr_80_io_en),
    .io_scan_mode(rvclkhdr_80_io_scan_mode)
  );
  rvclkhdr rvclkhdr_81 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_81_io_l1clk),
    .io_clk(rvclkhdr_81_io_clk),
    .io_en(rvclkhdr_81_io_en),
    .io_scan_mode(rvclkhdr_81_io_scan_mode)
  );
  rvclkhdr rvclkhdr_82 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_82_io_l1clk),
    .io_clk(rvclkhdr_82_io_clk),
    .io_en(rvclkhdr_82_io_en),
    .io_scan_mode(rvclkhdr_82_io_scan_mode)
  );
  rvclkhdr rvclkhdr_83 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_83_io_l1clk),
    .io_clk(rvclkhdr_83_io_clk),
    .io_en(rvclkhdr_83_io_en),
    .io_scan_mode(rvclkhdr_83_io_scan_mode)
  );
  rvclkhdr rvclkhdr_84 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_84_io_l1clk),
    .io_clk(rvclkhdr_84_io_clk),
    .io_en(rvclkhdr_84_io_en),
    .io_scan_mode(rvclkhdr_84_io_scan_mode)
  );
  rvclkhdr rvclkhdr_85 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_85_io_l1clk),
    .io_clk(rvclkhdr_85_io_clk),
    .io_en(rvclkhdr_85_io_en),
    .io_scan_mode(rvclkhdr_85_io_scan_mode)
  );
  rvclkhdr rvclkhdr_86 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_86_io_l1clk),
    .io_clk(rvclkhdr_86_io_clk),
    .io_en(rvclkhdr_86_io_en),
    .io_scan_mode(rvclkhdr_86_io_scan_mode)
  );
  rvclkhdr rvclkhdr_87 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_87_io_l1clk),
    .io_clk(rvclkhdr_87_io_clk),
    .io_en(rvclkhdr_87_io_en),
    .io_scan_mode(rvclkhdr_87_io_scan_mode)
  );
  rvclkhdr rvclkhdr_88 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_88_io_l1clk),
    .io_clk(rvclkhdr_88_io_clk),
    .io_en(rvclkhdr_88_io_en),
    .io_scan_mode(rvclkhdr_88_io_scan_mode)
  );
  rvclkhdr rvclkhdr_89 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_89_io_l1clk),
    .io_clk(rvclkhdr_89_io_clk),
    .io_en(rvclkhdr_89_io_en),
    .io_scan_mode(rvclkhdr_89_io_scan_mode)
  );
  rvclkhdr rvclkhdr_90 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_90_io_l1clk),
    .io_clk(rvclkhdr_90_io_clk),
    .io_en(rvclkhdr_90_io_en),
    .io_scan_mode(rvclkhdr_90_io_scan_mode)
  );
  rvclkhdr rvclkhdr_91 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_91_io_l1clk),
    .io_clk(rvclkhdr_91_io_clk),
    .io_en(rvclkhdr_91_io_en),
    .io_scan_mode(rvclkhdr_91_io_scan_mode)
  );
  rvclkhdr rvclkhdr_92 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_92_io_l1clk),
    .io_clk(rvclkhdr_92_io_clk),
    .io_en(rvclkhdr_92_io_en),
    .io_scan_mode(rvclkhdr_92_io_scan_mode)
  );
  rvclkhdr rvclkhdr_93 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_93_io_l1clk),
    .io_clk(rvclkhdr_93_io_clk),
    .io_en(rvclkhdr_93_io_en),
    .io_scan_mode(rvclkhdr_93_io_scan_mode)
  );
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 331:26]
  assign io_ifu_ic_mb_empty = _T_328 | _T_231; // @[el2_ifu_mem_ctl.scala 330:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 194:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3936; // @[el2_ifu_mem_ctl.scala 705:21]
  assign io_ifu_pmu_ic_miss = _T_9747; // @[el2_ifu_mem_ctl.scala 822:22]
  assign io_ifu_pmu_ic_hit = _T_9748; // @[el2_ifu_mem_ctl.scala 823:21]
  assign io_ifu_pmu_bus_error = _T_9749; // @[el2_ifu_mem_ctl.scala 824:24]
  assign io_ifu_pmu_bus_busy = _T_9753; // @[el2_ifu_mem_ctl.scala 825:23]
  assign io_ifu_pmu_bus_trxn = _T_9754; // @[el2_ifu_mem_ctl.scala 826:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 144:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 143:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 138:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 142:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 140:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 151:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 153:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 148:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 146:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 139:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 137:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 135:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 136:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 145:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 154:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 149:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 566:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2558; // @[el2_ifu_mem_ctl.scala 567:19]
  assign io_ifu_axi_araddr = _T_2560 & _T_2562; // @[el2_ifu_mem_ctl.scala 568:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 571:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 150:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 569:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 572:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 141:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 570:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 152:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 147:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 573:21]
  assign io_iccm_dma_ecc_error = iccm_dma_ecc_error; // @[el2_ifu_mem_ctl.scala 664:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 662:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 666:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 657:20]
  assign io_iccm_ready = _T_2656 & _T_2650; // @[el2_ifu_mem_ctl.scala 636:17]
  assign io_ic_rw_addr = _T_340 | _T_341; // @[el2_ifu_mem_ctl.scala 340:17]
  assign io_ic_wr_en = bus_ic_wr_en & _T_3922; // @[el2_ifu_mem_ctl.scala 704:15]
  assign io_ic_rd_en = _T_3914 | _T_3919; // @[el2_ifu_mem_ctl.scala 695:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 347:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 347:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 348:23]
  assign io_ifu_ic_debug_rd_data = _T_1211; // @[el2_ifu_mem_ctl.scala 356:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 829:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 831:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 832:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 830:25]
  assign io_ic_debug_way = _T_9766[1:0]; // @[el2_ifu_mem_ctl.scala 833:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_9740; // @[el2_ifu_mem_ctl.scala 817:19]
  assign io_iccm_rw_addr = _T_3060 ? io_dma_mem_addr[15:1] : _T_3067; // @[el2_ifu_mem_ctl.scala 668:19]
  assign io_iccm_wren = _T_2660 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 638:16]
  assign io_iccm_rden = _T_2664 | _T_2665; // @[el2_ifu_mem_ctl.scala 639:16]
  assign io_iccm_wr_data = _T_3042 ? _T_3043 : _T_3050; // @[el2_ifu_mem_ctl.scala 645:19]
  assign io_iccm_wr_size = _T_2670 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 641:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 291:15]
  assign io_ic_access_fault_f = _T_2443 & _T_319; // @[el2_ifu_mem_ctl.scala 388:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1273; // @[el2_ifu_mem_ctl.scala 389:29]
  assign io_iccm_rd_ecc_single_err = _T_3859 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 681:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 682:29]
  assign io_ic_error_start = _T_1199 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 350:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 193:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 192:24]
  assign io_ic_fetch_val_f = {_T_1281,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 392:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 385:16]
  assign io_ic_premux_data = ic_premux_data_temp[63:0]; // @[el2_ifu_mem_ctl.scala 382:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 383:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_9775; // @[el2_ifu_mem_ctl.scala 840:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2448; // @[el2_ifu_mem_ctl.scala 483:27]
  assign io_iccm_correction_state = _T_2476 ? 1'h0 : _GEN_43; // @[el2_ifu_mem_ctl.scala 518:28 el2_ifu_mem_ctl.scala 531:32 el2_ifu_mem_ctl.scala 538:32 el2_ifu_mem_ctl.scala 545:32]
  assign rvclkhdr_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_io_en = ic_debug_rd_en_ff; // @[el2_lib.scala 485:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_1_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_1_io_en = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_lib.scala 485:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_2_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_2_io_en = _T_2 | scnd_miss_req; // @[el2_lib.scala 485:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_3_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_3_io_en = _T_309 | io_dec_tlu_force_halt; // @[el2_lib.scala 485:16]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_4_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_4_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_5_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_5_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_6_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_6_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_7_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_7_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_8_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_8_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_9_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_9_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_10_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_10_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_11_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_11_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_12_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_12_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_13_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_13_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_14_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_14_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_15_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_15_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_16_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_16_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_17_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_17_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_18_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_18_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_19_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_19_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_20_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_20_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_21_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_21_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_22_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_22_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_23_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_23_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_24_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_24_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_25_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_25_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_26_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_26_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_26_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_27_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_27_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_27_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_28_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_28_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_28_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_29_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_29_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_29_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_30_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_30_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_30_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_31_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_31_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_31_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_32_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_32_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_32_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_33_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_33_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_33_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_34_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_34_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_34_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_35_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_35_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_35_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_36_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_36_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_36_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_37_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_37_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_37_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_38_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_38_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_38_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_39_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_39_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_39_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_40_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_40_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_40_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_41_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_41_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_41_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_42_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_42_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_42_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_43_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_43_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_43_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_44_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_44_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_44_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_45_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_45_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_45_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_46_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_46_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_46_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_47_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_47_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_47_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_48_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_48_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_48_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_49_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_49_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_49_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_50_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_50_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_50_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_51_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_51_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_51_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_52_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_52_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_52_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_53_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_53_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_53_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_54_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_54_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_54_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_55_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_55_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_55_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_56_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_56_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_56_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_57_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_57_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_57_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_58_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_58_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_58_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_59_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_59_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_59_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_60_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_60_io_en = bus_ifu_wr_en & _T_1284; // @[el2_lib.scala 485:16]
  assign rvclkhdr_60_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_61_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_61_io_en = bus_ifu_wr_en & _T_1285; // @[el2_lib.scala 485:16]
  assign rvclkhdr_61_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_62_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_62_io_en = bus_ifu_wr_en & _T_1286; // @[el2_lib.scala 485:16]
  assign rvclkhdr_62_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_63_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_63_io_en = bus_ifu_wr_en & _T_1287; // @[el2_lib.scala 485:16]
  assign rvclkhdr_63_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_64_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_64_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_64_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_65_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_65_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_65_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_66_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_66_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_66_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_67_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_67_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_67_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_68_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_68_io_en = io_ifu_bus_clk_en; // @[el2_lib.scala 485:16]
  assign rvclkhdr_68_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_69_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_69_io_en = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_lib.scala 485:16]
  assign rvclkhdr_69_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_70_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_70_io_en = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_lib.scala 485:16]
  assign rvclkhdr_70_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_71_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_71_io_en = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_lib.scala 485:16]
  assign rvclkhdr_71_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_72_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_72_io_en = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_lib.scala 485:16]
  assign rvclkhdr_72_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_73_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_73_io_en = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_lib.scala 485:16]
  assign rvclkhdr_73_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_74_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_74_io_en = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_lib.scala 485:16]
  assign rvclkhdr_74_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_75_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_75_io_en = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_lib.scala 485:16]
  assign rvclkhdr_75_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_76_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_76_io_en = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_lib.scala 485:16]
  assign rvclkhdr_76_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_77_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_77_io_en = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_lib.scala 485:16]
  assign rvclkhdr_77_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_78_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_78_io_en = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_lib.scala 485:16]
  assign rvclkhdr_78_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_79_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_79_io_en = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_lib.scala 485:16]
  assign rvclkhdr_79_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_80_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_80_io_en = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_lib.scala 485:16]
  assign rvclkhdr_80_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_81_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_81_io_en = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_lib.scala 485:16]
  assign rvclkhdr_81_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_82_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_82_io_en = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_lib.scala 485:16]
  assign rvclkhdr_82_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_83_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_83_io_en = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_lib.scala 485:16]
  assign rvclkhdr_83_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_84_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_84_io_en = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_lib.scala 485:16]
  assign rvclkhdr_84_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_85_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_85_io_en = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_lib.scala 485:16]
  assign rvclkhdr_85_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_86_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_86_io_en = tag_valid_clken_0[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_86_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_87_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_87_io_en = tag_valid_clken_0[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_87_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_88_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_88_io_en = tag_valid_clken_1[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_88_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_89_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_89_io_en = tag_valid_clken_1[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_89_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_90_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_90_io_en = tag_valid_clken_2[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_90_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_91_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_91_io_en = tag_valid_clken_2[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_91_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_92_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_92_io_en = tag_valid_clken_3[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_92_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_93_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_93_io_en = tag_valid_clken_3[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_93_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ifu_ic_rw_int_addr_ff = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  way_status_out_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_status_out_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_status_out_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_status_out_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_status_out_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_status_out_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_status_out_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_status_out_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_status_out_8 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_status_out_9 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_status_out_10 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_status_out_11 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_status_out_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_status_out_13 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_status_out_14 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_status_out_15 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_status_out_16 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_status_out_17 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_status_out_18 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_status_out_19 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_status_out_20 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_status_out_21 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_status_out_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_status_out_23 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_status_out_24 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_status_out_25 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_status_out_26 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_status_out_27 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_status_out_28 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_status_out_29 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_status_out_30 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_status_out_31 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_status_out_32 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_status_out_33 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_status_out_34 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_status_out_35 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_status_out_36 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_status_out_37 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_status_out_38 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_status_out_39 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_status_out_40 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_status_out_41 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way_status_out_42 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way_status_out_43 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way_status_out_44 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way_status_out_45 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way_status_out_46 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way_status_out_47 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way_status_out_48 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way_status_out_49 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way_status_out_50 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way_status_out_51 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way_status_out_52 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way_status_out_53 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way_status_out_54 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way_status_out_55 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way_status_out_56 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way_status_out_57 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way_status_out_58 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way_status_out_59 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way_status_out_60 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way_status_out_61 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way_status_out_62 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way_status_out_63 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way_status_out_64 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way_status_out_65 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way_status_out_66 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way_status_out_67 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way_status_out_68 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way_status_out_69 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way_status_out_70 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way_status_out_71 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way_status_out_72 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way_status_out_73 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way_status_out_74 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way_status_out_75 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way_status_out_76 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way_status_out_77 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way_status_out_78 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way_status_out_79 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way_status_out_80 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way_status_out_81 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way_status_out_82 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way_status_out_83 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way_status_out_84 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way_status_out_85 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way_status_out_86 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way_status_out_87 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way_status_out_88 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way_status_out_89 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way_status_out_90 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way_status_out_91 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way_status_out_92 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way_status_out_93 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way_status_out_94 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way_status_out_95 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way_status_out_96 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way_status_out_97 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way_status_out_98 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way_status_out_99 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way_status_out_100 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way_status_out_101 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way_status_out_102 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way_status_out_103 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way_status_out_104 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way_status_out_105 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way_status_out_106 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way_status_out_107 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  way_status_out_108 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  way_status_out_109 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way_status_out_110 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way_status_out_111 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way_status_out_112 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way_status_out_113 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way_status_out_114 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way_status_out_115 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way_status_out_116 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way_status_out_117 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way_status_out_118 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way_status_out_119 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way_status_out_120 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way_status_out_121 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way_status_out_122 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way_status_out_123 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way_status_out_124 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way_status_out_125 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way_status_out_126 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way_status_out_127 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  tagv_mb_scnd_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_152[30:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  reset_ic_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  miss_addr = _RAND_160[25:0];
  _RAND_161 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_163[0:0];
  _RAND_164 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_164[63:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_441[0:0];
  _RAND_442 = {3{`RANDOM}};
  _T_1211 = _RAND_442[70:0];
  _RAND_443 = {1{`RANDOM}};
  ifc_region_acc_fault_memory_f = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_444[6:0];
  _RAND_445 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  bus_cmd_req_hold = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_448[2:0];
  _RAND_449 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_451[0:0];
  _RAND_452 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_452[38:0];
  _RAND_453 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_454[2:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_dma_rtag_temp = _RAND_455[2:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_dma_rvalid_temp = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_dma_ecc_error = _RAND_457[0:0];
  _RAND_458 = {2{`RANDOM}};
  iccm_dma_rdata_temp = _RAND_458[63:0];
  _RAND_459 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_459[13:0];
  _RAND_460 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_461[13:0];
  _RAND_462 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_462[6:0];
  _RAND_463 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  way_status_new_ff = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  ic_valid_ff = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_9747 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_9748 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_9749 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  _T_9753 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  _T_9754 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  _T_9775 = _RAND_472[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    flush_final_f = 1'h0;
  end
  if (reset) begin
    ifc_fetch_req_f_raw = 1'h0;
  end
  if (reset) begin
    miss_state = 3'h0;
  end
  if (reset) begin
    scnd_miss_req_q = 1'h0;
  end
  if (reset) begin
    ifu_fetch_addr_int_f = 31'h0;
  end
  if (reset) begin
    ifc_iccm_access_f = 1'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_in = 1'h0;
  end
  if (reset) begin
    dma_iccm_req_f = 1'h0;
  end
  if (reset) begin
    perr_state = 3'h0;
  end
  if (reset) begin
    err_stop_state = 2'h0;
  end
  if (reset) begin
    reset_all_tags = 1'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_final_f = 1'h0;
  end
  if (reset) begin
    ifu_bus_rvalid_unq_ff = 1'h0;
  end
  if (reset) begin
    bus_ifu_bus_clk_en_ff = 1'h0;
  end
  if (reset) begin
    uncacheable_miss_ff = 1'h0;
  end
  if (reset) begin
    bus_data_beat_count = 3'h0;
  end
  if (reset) begin
    ic_miss_buff_data_valid = 8'h0;
  end
  if (reset) begin
    last_data_recieved_ff = 1'h0;
  end
  if (reset) begin
    sel_mb_addr_ff = 1'h0;
  end
  if (reset) begin
    way_status_mb_scnd_ff = 1'h0;
  end
  if (reset) begin
    ifu_ic_rw_int_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_out_0 = 1'h0;
  end
  if (reset) begin
    way_status_out_1 = 1'h0;
  end
  if (reset) begin
    way_status_out_2 = 1'h0;
  end
  if (reset) begin
    way_status_out_3 = 1'h0;
  end
  if (reset) begin
    way_status_out_4 = 1'h0;
  end
  if (reset) begin
    way_status_out_5 = 1'h0;
  end
  if (reset) begin
    way_status_out_6 = 1'h0;
  end
  if (reset) begin
    way_status_out_7 = 1'h0;
  end
  if (reset) begin
    way_status_out_8 = 1'h0;
  end
  if (reset) begin
    way_status_out_9 = 1'h0;
  end
  if (reset) begin
    way_status_out_10 = 1'h0;
  end
  if (reset) begin
    way_status_out_11 = 1'h0;
  end
  if (reset) begin
    way_status_out_12 = 1'h0;
  end
  if (reset) begin
    way_status_out_13 = 1'h0;
  end
  if (reset) begin
    way_status_out_14 = 1'h0;
  end
  if (reset) begin
    way_status_out_15 = 1'h0;
  end
  if (reset) begin
    way_status_out_16 = 1'h0;
  end
  if (reset) begin
    way_status_out_17 = 1'h0;
  end
  if (reset) begin
    way_status_out_18 = 1'h0;
  end
  if (reset) begin
    way_status_out_19 = 1'h0;
  end
  if (reset) begin
    way_status_out_20 = 1'h0;
  end
  if (reset) begin
    way_status_out_21 = 1'h0;
  end
  if (reset) begin
    way_status_out_22 = 1'h0;
  end
  if (reset) begin
    way_status_out_23 = 1'h0;
  end
  if (reset) begin
    way_status_out_24 = 1'h0;
  end
  if (reset) begin
    way_status_out_25 = 1'h0;
  end
  if (reset) begin
    way_status_out_26 = 1'h0;
  end
  if (reset) begin
    way_status_out_27 = 1'h0;
  end
  if (reset) begin
    way_status_out_28 = 1'h0;
  end
  if (reset) begin
    way_status_out_29 = 1'h0;
  end
  if (reset) begin
    way_status_out_30 = 1'h0;
  end
  if (reset) begin
    way_status_out_31 = 1'h0;
  end
  if (reset) begin
    way_status_out_32 = 1'h0;
  end
  if (reset) begin
    way_status_out_33 = 1'h0;
  end
  if (reset) begin
    way_status_out_34 = 1'h0;
  end
  if (reset) begin
    way_status_out_35 = 1'h0;
  end
  if (reset) begin
    way_status_out_36 = 1'h0;
  end
  if (reset) begin
    way_status_out_37 = 1'h0;
  end
  if (reset) begin
    way_status_out_38 = 1'h0;
  end
  if (reset) begin
    way_status_out_39 = 1'h0;
  end
  if (reset) begin
    way_status_out_40 = 1'h0;
  end
  if (reset) begin
    way_status_out_41 = 1'h0;
  end
  if (reset) begin
    way_status_out_42 = 1'h0;
  end
  if (reset) begin
    way_status_out_43 = 1'h0;
  end
  if (reset) begin
    way_status_out_44 = 1'h0;
  end
  if (reset) begin
    way_status_out_45 = 1'h0;
  end
  if (reset) begin
    way_status_out_46 = 1'h0;
  end
  if (reset) begin
    way_status_out_47 = 1'h0;
  end
  if (reset) begin
    way_status_out_48 = 1'h0;
  end
  if (reset) begin
    way_status_out_49 = 1'h0;
  end
  if (reset) begin
    way_status_out_50 = 1'h0;
  end
  if (reset) begin
    way_status_out_51 = 1'h0;
  end
  if (reset) begin
    way_status_out_52 = 1'h0;
  end
  if (reset) begin
    way_status_out_53 = 1'h0;
  end
  if (reset) begin
    way_status_out_54 = 1'h0;
  end
  if (reset) begin
    way_status_out_55 = 1'h0;
  end
  if (reset) begin
    way_status_out_56 = 1'h0;
  end
  if (reset) begin
    way_status_out_57 = 1'h0;
  end
  if (reset) begin
    way_status_out_58 = 1'h0;
  end
  if (reset) begin
    way_status_out_59 = 1'h0;
  end
  if (reset) begin
    way_status_out_60 = 1'h0;
  end
  if (reset) begin
    way_status_out_61 = 1'h0;
  end
  if (reset) begin
    way_status_out_62 = 1'h0;
  end
  if (reset) begin
    way_status_out_63 = 1'h0;
  end
  if (reset) begin
    way_status_out_64 = 1'h0;
  end
  if (reset) begin
    way_status_out_65 = 1'h0;
  end
  if (reset) begin
    way_status_out_66 = 1'h0;
  end
  if (reset) begin
    way_status_out_67 = 1'h0;
  end
  if (reset) begin
    way_status_out_68 = 1'h0;
  end
  if (reset) begin
    way_status_out_69 = 1'h0;
  end
  if (reset) begin
    way_status_out_70 = 1'h0;
  end
  if (reset) begin
    way_status_out_71 = 1'h0;
  end
  if (reset) begin
    way_status_out_72 = 1'h0;
  end
  if (reset) begin
    way_status_out_73 = 1'h0;
  end
  if (reset) begin
    way_status_out_74 = 1'h0;
  end
  if (reset) begin
    way_status_out_75 = 1'h0;
  end
  if (reset) begin
    way_status_out_76 = 1'h0;
  end
  if (reset) begin
    way_status_out_77 = 1'h0;
  end
  if (reset) begin
    way_status_out_78 = 1'h0;
  end
  if (reset) begin
    way_status_out_79 = 1'h0;
  end
  if (reset) begin
    way_status_out_80 = 1'h0;
  end
  if (reset) begin
    way_status_out_81 = 1'h0;
  end
  if (reset) begin
    way_status_out_82 = 1'h0;
  end
  if (reset) begin
    way_status_out_83 = 1'h0;
  end
  if (reset) begin
    way_status_out_84 = 1'h0;
  end
  if (reset) begin
    way_status_out_85 = 1'h0;
  end
  if (reset) begin
    way_status_out_86 = 1'h0;
  end
  if (reset) begin
    way_status_out_87 = 1'h0;
  end
  if (reset) begin
    way_status_out_88 = 1'h0;
  end
  if (reset) begin
    way_status_out_89 = 1'h0;
  end
  if (reset) begin
    way_status_out_90 = 1'h0;
  end
  if (reset) begin
    way_status_out_91 = 1'h0;
  end
  if (reset) begin
    way_status_out_92 = 1'h0;
  end
  if (reset) begin
    way_status_out_93 = 1'h0;
  end
  if (reset) begin
    way_status_out_94 = 1'h0;
  end
  if (reset) begin
    way_status_out_95 = 1'h0;
  end
  if (reset) begin
    way_status_out_96 = 1'h0;
  end
  if (reset) begin
    way_status_out_97 = 1'h0;
  end
  if (reset) begin
    way_status_out_98 = 1'h0;
  end
  if (reset) begin
    way_status_out_99 = 1'h0;
  end
  if (reset) begin
    way_status_out_100 = 1'h0;
  end
  if (reset) begin
    way_status_out_101 = 1'h0;
  end
  if (reset) begin
    way_status_out_102 = 1'h0;
  end
  if (reset) begin
    way_status_out_103 = 1'h0;
  end
  if (reset) begin
    way_status_out_104 = 1'h0;
  end
  if (reset) begin
    way_status_out_105 = 1'h0;
  end
  if (reset) begin
    way_status_out_106 = 1'h0;
  end
  if (reset) begin
    way_status_out_107 = 1'h0;
  end
  if (reset) begin
    way_status_out_108 = 1'h0;
  end
  if (reset) begin
    way_status_out_109 = 1'h0;
  end
  if (reset) begin
    way_status_out_110 = 1'h0;
  end
  if (reset) begin
    way_status_out_111 = 1'h0;
  end
  if (reset) begin
    way_status_out_112 = 1'h0;
  end
  if (reset) begin
    way_status_out_113 = 1'h0;
  end
  if (reset) begin
    way_status_out_114 = 1'h0;
  end
  if (reset) begin
    way_status_out_115 = 1'h0;
  end
  if (reset) begin
    way_status_out_116 = 1'h0;
  end
  if (reset) begin
    way_status_out_117 = 1'h0;
  end
  if (reset) begin
    way_status_out_118 = 1'h0;
  end
  if (reset) begin
    way_status_out_119 = 1'h0;
  end
  if (reset) begin
    way_status_out_120 = 1'h0;
  end
  if (reset) begin
    way_status_out_121 = 1'h0;
  end
  if (reset) begin
    way_status_out_122 = 1'h0;
  end
  if (reset) begin
    way_status_out_123 = 1'h0;
  end
  if (reset) begin
    way_status_out_124 = 1'h0;
  end
  if (reset) begin
    way_status_out_125 = 1'h0;
  end
  if (reset) begin
    way_status_out_126 = 1'h0;
  end
  if (reset) begin
    way_status_out_127 = 1'h0;
  end
  if (reset) begin
    tagv_mb_scnd_ff = 2'h0;
  end
  if (reset) begin
    uncacheable_miss_scnd_ff = 1'h0;
  end
  if (reset) begin
    imb_scnd_ff = 31'h0;
  end
  if (reset) begin
    ifu_bus_rid_ff = 3'h0;
  end
  if (reset) begin
    ifu_bus_rresp_ff = 2'h0;
  end
  if (reset) begin
    ifu_wr_data_comb_err_ff = 1'h0;
  end
  if (reset) begin
    way_status_mb_ff = 1'h0;
  end
  if (reset) begin
    tagv_mb_ff = 2'h0;
  end
  if (reset) begin
    fetch_uncacheable_ff = 1'h0;
  end
  if (reset) begin
    miss_addr = 26'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_f = 1'h0;
  end
  if (reset) begin
    bus_rd_addr_count = 3'h0;
  end
  if (reset) begin
    ic_act_miss_f_delayed = 1'h0;
  end
  if (reset) begin
    ifu_bus_rdata_ff = 64'h0;
  end
  if (reset) begin
    ic_miss_buff_data_0 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_1 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_2 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_3 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_4 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_5 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_6 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_7 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_8 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_9 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_10 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_11 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_12 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_13 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_14 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_15 = 32'h0;
  end
  if (reset) begin
    ic_crit_wd_rdy_new_ff = 1'h0;
  end
  if (reset) begin
    ic_miss_buff_data_error = 8'h0;
  end
  if (reset) begin
    ic_debug_ict_array_sel_ff = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_127 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_127 = 1'h0;
  end
  if (reset) begin
    ic_debug_way_ff = 2'h0;
  end
  if (reset) begin
    ic_debug_rd_en_ff = 1'h0;
  end
  if (reset) begin
    _T_1211 = 71'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_memory_f = 1'h0;
  end
  if (reset) begin
    perr_ic_index_ff = 7'h0;
  end
  if (reset) begin
    dma_sb_err_state_ff = 1'h0;
  end
  if (reset) begin
    bus_cmd_req_hold = 1'h0;
  end
  if (reset) begin
    ifu_bus_cmd_valid = 1'h0;
  end
  if (reset) begin
    bus_cmd_beat_count = 3'h0;
  end
  if (reset) begin
    ifu_bus_arready_unq_ff = 1'h0;
  end
  if (reset) begin
    ifu_bus_arvalid_ff = 1'h0;
  end
  if (reset) begin
    ifc_dma_access_ok_prev = 1'h0;
  end
  if (reset) begin
    iccm_ecc_corr_data_ff = 39'h0;
  end
  if (reset) begin
    dma_mem_addr_ff = 2'h0;
  end
  if (reset) begin
    dma_mem_tag_ff = 3'h0;
  end
  if (reset) begin
    iccm_dma_rtag_temp = 3'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_temp = 1'h0;
  end
  if (reset) begin
    iccm_dma_ecc_error = 1'h0;
  end
  if (reset) begin
    iccm_dma_rdata_temp = 64'h0;
  end
  if (reset) begin
    iccm_ecc_corr_index_ff = 14'h0;
  end
  if (reset) begin
    iccm_rd_ecc_single_err_ff = 1'h0;
  end
  if (reset) begin
    iccm_rw_addr_f = 14'h0;
  end
  if (reset) begin
    ifu_status_wr_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_wr_en_ff = 1'h0;
  end
  if (reset) begin
    way_status_new_ff = 1'h0;
  end
  if (reset) begin
    ifu_tag_wren_ff = 2'h0;
  end
  if (reset) begin
    ic_valid_ff = 1'h0;
  end
  if (reset) begin
    _T_9747 = 1'h0;
  end
  if (reset) begin
    _T_9748 = 1'h0;
  end
  if (reset) begin
    _T_9749 = 1'h0;
  end
  if (reset) begin
    _T_9753 = 1'h0;
  end
  if (reset) begin
    _T_9754 = 1'h0;
  end
  if (reset) begin
    _T_9775 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge rvclkhdr_2_io_l1clk) begin
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge clock) begin
    reset_ic_ff <= _T_298 & _T_299;
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= _T_317 & _T_318;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= _T_22 & _T_319;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2659 & _T_2663;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2451) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2453) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2463) begin
        perr_state <= 3'h0;
      end else if (_T_2466) begin
        if (_T_2468) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2472) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2476) begin
        err_stop_state <= 2'h1;
      end else if (_T_2481) begin
        if (_T_2483) begin
          err_stop_state <= 2'h0;
        end else if (_T_2504) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2508) begin
        if (_T_2483) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2525) begin
        if (_T_2529) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf | ifc_region_acc_fault_memory_bf;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= _T_2581 | _T_2582;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= {_T_1353,ic_miss_buff_data_valid_in_0};
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= _T_2589 | _T_2591;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= _T_334 | reset_tag_valid_for_miss;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_ic_rw_int_addr_ff <= 7'h0;
    end else if (_T_3945) begin
      ifu_ic_rw_int_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_ic_rw_int_addr_ff <= ifu_ic_rw_int_addr[11:5];
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_0 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_0 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_1 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_1 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_2 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_2 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_3 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_3 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_4 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_4 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_5 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_5 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_6 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_6 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_7 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_7 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_8 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_8 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_9 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_9 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_10 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_10 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_11 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_11 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_12 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_12 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_13 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_13 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_14 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_14 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_15 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_15 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_16 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_16 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_17 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_17 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_18 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_18 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_19 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_19 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_20 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_20 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_21 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_21 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_22 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_22 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_23 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_23 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_24 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_24 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_25 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_25 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_26 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_26 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_27 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_27 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_28 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_28 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_29 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_29 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_30 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_30 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_31 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_31 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_32 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_32 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_33 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_33 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_34 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_34 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_35 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_35 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_36 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_36 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_37 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_37 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_38 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_38 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_39 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_39 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_40 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_40 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_41 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_41 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_42 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_42 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_43 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_43 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_44 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_44 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_45 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_45 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_46 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_46 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_47 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_47 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_48 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_48 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_49 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_49 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_50 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_50 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_51 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_51 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_52 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_52 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_53 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_53 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_54 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_54 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_55 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_55 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_56 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_56 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_57 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_57 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_58 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_58 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_59 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_59 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_60 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_60 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_61 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_61 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_62 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_62 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_63 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_63 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_64 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_64 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_65 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_65 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_66 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_66 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_67 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_67 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_68 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_68 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_69 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_69 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_70 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_70 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_71 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_71 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_72 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_72 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_73 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_73 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_74 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_74 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_75 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_75 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_76 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_76 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_77 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_77 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_78 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_78 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_79 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_79 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_80 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_80 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_81 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_81 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_82 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_82 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_83 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_83 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_84 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_84 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_85 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_85 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_86 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_86 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_87 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_87 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_88 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_88 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_89 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_89 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_90 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_90 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_91 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_91 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_92 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_92 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_93 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_93 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_94 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_94 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_95 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_95 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_96 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_96 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_97 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_97 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_98 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_98 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_99 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_99 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_100 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_100 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_101 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_101 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_102 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_102 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_103 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_103 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_104 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_104 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_105 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_105 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_106 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_106 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_107 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_107 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_108 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_108 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_109 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_109 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_110 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_110 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_111 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_111 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_112 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_112 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_113 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_113 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_114 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_114 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_115 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_115 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_116 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_116 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_117 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_117 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_118 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_118 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_119 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_119 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_120 <= 1'h0;
    end else if (_T_3969) begin
      way_status_out_120 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_121 <= 1'h0;
    end else if (_T_3973) begin
      way_status_out_121 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_122 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_122 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_123 <= 1'h0;
    end else if (_T_3981) begin
      way_status_out_123 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_124 <= 1'h0;
    end else if (_T_3985) begin
      way_status_out_124 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_125 <= 1'h0;
    end else if (_T_3989) begin
      way_status_out_125 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_126 <= 1'h0;
    end else if (_T_3993) begin
      way_status_out_126 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_127 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_127 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      tagv_mb_scnd_ff <= 2'h0;
    end else if (!(_T_19)) begin
      tagv_mb_scnd_ff <= _T_198;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err_data & _T_2577;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_290;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= _T_295;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_231) begin
      bus_rd_addr_count <= imb_ff[4:2];
    end else if (scnd_miss_req_q) begin
      bus_rd_addr_count <= imb_scnd_ff[4:2];
    end else if (bus_cmd_sent) begin
      bus_rd_addr_count <= _T_2597;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= _T_233 & _T_209;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_40_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_40_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_49_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_49_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_58_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_58_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_67_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_67_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= _T_1509 | _T_1514;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= {_T_1393,ic_miss_buff_data_error_in_0};
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else begin
      ic_debug_ict_array_sel_ff <= io_ic_debug_rd_en & io_ic_debug_tag_array;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5590) begin
      ic_tag_valid_out_1_0 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5605) begin
      ic_tag_valid_out_1_1 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5620) begin
      ic_tag_valid_out_1_2 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5635) begin
      ic_tag_valid_out_1_3 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5650) begin
      ic_tag_valid_out_1_4 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5665) begin
      ic_tag_valid_out_1_5 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5680) begin
      ic_tag_valid_out_1_6 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5695) begin
      ic_tag_valid_out_1_7 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5710) begin
      ic_tag_valid_out_1_8 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5725) begin
      ic_tag_valid_out_1_9 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5740) begin
      ic_tag_valid_out_1_10 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5755) begin
      ic_tag_valid_out_1_11 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5770) begin
      ic_tag_valid_out_1_12 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5785) begin
      ic_tag_valid_out_1_13 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5800) begin
      ic_tag_valid_out_1_14 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5815) begin
      ic_tag_valid_out_1_15 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5830) begin
      ic_tag_valid_out_1_16 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5845) begin
      ic_tag_valid_out_1_17 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5860) begin
      ic_tag_valid_out_1_18 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5875) begin
      ic_tag_valid_out_1_19 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5890) begin
      ic_tag_valid_out_1_20 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5905) begin
      ic_tag_valid_out_1_21 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5920) begin
      ic_tag_valid_out_1_22 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5935) begin
      ic_tag_valid_out_1_23 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_5950) begin
      ic_tag_valid_out_1_24 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_5965) begin
      ic_tag_valid_out_1_25 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_5980) begin
      ic_tag_valid_out_1_26 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_5995) begin
      ic_tag_valid_out_1_27 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6010) begin
      ic_tag_valid_out_1_28 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6025) begin
      ic_tag_valid_out_1_29 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6040) begin
      ic_tag_valid_out_1_30 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6055) begin
      ic_tag_valid_out_1_31 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6550) begin
      ic_tag_valid_out_1_32 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6565) begin
      ic_tag_valid_out_1_33 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6580) begin
      ic_tag_valid_out_1_34 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6595) begin
      ic_tag_valid_out_1_35 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6610) begin
      ic_tag_valid_out_1_36 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6625) begin
      ic_tag_valid_out_1_37 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6640) begin
      ic_tag_valid_out_1_38 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6655) begin
      ic_tag_valid_out_1_39 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6670) begin
      ic_tag_valid_out_1_40 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6685) begin
      ic_tag_valid_out_1_41 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6700) begin
      ic_tag_valid_out_1_42 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6715) begin
      ic_tag_valid_out_1_43 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6730) begin
      ic_tag_valid_out_1_44 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6745) begin
      ic_tag_valid_out_1_45 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6760) begin
      ic_tag_valid_out_1_46 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6775) begin
      ic_tag_valid_out_1_47 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6790) begin
      ic_tag_valid_out_1_48 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6805) begin
      ic_tag_valid_out_1_49 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6820) begin
      ic_tag_valid_out_1_50 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6835) begin
      ic_tag_valid_out_1_51 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6850) begin
      ic_tag_valid_out_1_52 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6865) begin
      ic_tag_valid_out_1_53 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6880) begin
      ic_tag_valid_out_1_54 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6895) begin
      ic_tag_valid_out_1_55 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6910) begin
      ic_tag_valid_out_1_56 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6925) begin
      ic_tag_valid_out_1_57 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6940) begin
      ic_tag_valid_out_1_58 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_6955) begin
      ic_tag_valid_out_1_59 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_6970) begin
      ic_tag_valid_out_1_60 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_6985) begin
      ic_tag_valid_out_1_61 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7000) begin
      ic_tag_valid_out_1_62 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7015) begin
      ic_tag_valid_out_1_63 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7510) begin
      ic_tag_valid_out_1_64 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7525) begin
      ic_tag_valid_out_1_65 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7540) begin
      ic_tag_valid_out_1_66 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7555) begin
      ic_tag_valid_out_1_67 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7570) begin
      ic_tag_valid_out_1_68 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7585) begin
      ic_tag_valid_out_1_69 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7600) begin
      ic_tag_valid_out_1_70 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7615) begin
      ic_tag_valid_out_1_71 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7630) begin
      ic_tag_valid_out_1_72 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7645) begin
      ic_tag_valid_out_1_73 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7660) begin
      ic_tag_valid_out_1_74 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7675) begin
      ic_tag_valid_out_1_75 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7690) begin
      ic_tag_valid_out_1_76 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7705) begin
      ic_tag_valid_out_1_77 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7720) begin
      ic_tag_valid_out_1_78 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7735) begin
      ic_tag_valid_out_1_79 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7750) begin
      ic_tag_valid_out_1_80 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7765) begin
      ic_tag_valid_out_1_81 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7780) begin
      ic_tag_valid_out_1_82 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7795) begin
      ic_tag_valid_out_1_83 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7810) begin
      ic_tag_valid_out_1_84 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7825) begin
      ic_tag_valid_out_1_85 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7840) begin
      ic_tag_valid_out_1_86 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7855) begin
      ic_tag_valid_out_1_87 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_7870) begin
      ic_tag_valid_out_1_88 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_7885) begin
      ic_tag_valid_out_1_89 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_7900) begin
      ic_tag_valid_out_1_90 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_7915) begin
      ic_tag_valid_out_1_91 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_7930) begin
      ic_tag_valid_out_1_92 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_7945) begin
      ic_tag_valid_out_1_93 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_7960) begin
      ic_tag_valid_out_1_94 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_7975) begin
      ic_tag_valid_out_1_95 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8470) begin
      ic_tag_valid_out_1_96 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8485) begin
      ic_tag_valid_out_1_97 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8500) begin
      ic_tag_valid_out_1_98 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8515) begin
      ic_tag_valid_out_1_99 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8530) begin
      ic_tag_valid_out_1_100 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8545) begin
      ic_tag_valid_out_1_101 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8560) begin
      ic_tag_valid_out_1_102 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8575) begin
      ic_tag_valid_out_1_103 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8590) begin
      ic_tag_valid_out_1_104 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8605) begin
      ic_tag_valid_out_1_105 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8620) begin
      ic_tag_valid_out_1_106 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8635) begin
      ic_tag_valid_out_1_107 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8650) begin
      ic_tag_valid_out_1_108 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8665) begin
      ic_tag_valid_out_1_109 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8680) begin
      ic_tag_valid_out_1_110 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8695) begin
      ic_tag_valid_out_1_111 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8710) begin
      ic_tag_valid_out_1_112 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8725) begin
      ic_tag_valid_out_1_113 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8740) begin
      ic_tag_valid_out_1_114 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_8755) begin
      ic_tag_valid_out_1_115 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_8770) begin
      ic_tag_valid_out_1_116 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_8785) begin
      ic_tag_valid_out_1_117 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_8800) begin
      ic_tag_valid_out_1_118 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_8815) begin
      ic_tag_valid_out_1_119 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_8830) begin
      ic_tag_valid_out_1_120 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_8845) begin
      ic_tag_valid_out_1_121 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_8860) begin
      ic_tag_valid_out_1_122 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_8875) begin
      ic_tag_valid_out_1_123 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_8890) begin
      ic_tag_valid_out_1_124 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_8905) begin
      ic_tag_valid_out_1_125 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_8920) begin
      ic_tag_valid_out_1_126 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_8935) begin
      ic_tag_valid_out_1_127 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5110) begin
      ic_tag_valid_out_0_0 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5125) begin
      ic_tag_valid_out_0_1 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5140) begin
      ic_tag_valid_out_0_2 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5155) begin
      ic_tag_valid_out_0_3 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5170) begin
      ic_tag_valid_out_0_4 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5185) begin
      ic_tag_valid_out_0_5 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5200) begin
      ic_tag_valid_out_0_6 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5215) begin
      ic_tag_valid_out_0_7 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5230) begin
      ic_tag_valid_out_0_8 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5245) begin
      ic_tag_valid_out_0_9 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5260) begin
      ic_tag_valid_out_0_10 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5275) begin
      ic_tag_valid_out_0_11 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5290) begin
      ic_tag_valid_out_0_12 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5305) begin
      ic_tag_valid_out_0_13 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5320) begin
      ic_tag_valid_out_0_14 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5335) begin
      ic_tag_valid_out_0_15 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5350) begin
      ic_tag_valid_out_0_16 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5365) begin
      ic_tag_valid_out_0_17 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5380) begin
      ic_tag_valid_out_0_18 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5395) begin
      ic_tag_valid_out_0_19 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5410) begin
      ic_tag_valid_out_0_20 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5425) begin
      ic_tag_valid_out_0_21 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5440) begin
      ic_tag_valid_out_0_22 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5455) begin
      ic_tag_valid_out_0_23 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5470) begin
      ic_tag_valid_out_0_24 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5485) begin
      ic_tag_valid_out_0_25 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5500) begin
      ic_tag_valid_out_0_26 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5515) begin
      ic_tag_valid_out_0_27 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5530) begin
      ic_tag_valid_out_0_28 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5545) begin
      ic_tag_valid_out_0_29 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5560) begin
      ic_tag_valid_out_0_30 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5575) begin
      ic_tag_valid_out_0_31 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6070) begin
      ic_tag_valid_out_0_32 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6085) begin
      ic_tag_valid_out_0_33 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6100) begin
      ic_tag_valid_out_0_34 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6115) begin
      ic_tag_valid_out_0_35 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6130) begin
      ic_tag_valid_out_0_36 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6145) begin
      ic_tag_valid_out_0_37 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6160) begin
      ic_tag_valid_out_0_38 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6175) begin
      ic_tag_valid_out_0_39 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6190) begin
      ic_tag_valid_out_0_40 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6205) begin
      ic_tag_valid_out_0_41 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6220) begin
      ic_tag_valid_out_0_42 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6235) begin
      ic_tag_valid_out_0_43 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6250) begin
      ic_tag_valid_out_0_44 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6265) begin
      ic_tag_valid_out_0_45 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6280) begin
      ic_tag_valid_out_0_46 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6295) begin
      ic_tag_valid_out_0_47 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6310) begin
      ic_tag_valid_out_0_48 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6325) begin
      ic_tag_valid_out_0_49 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6340) begin
      ic_tag_valid_out_0_50 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6355) begin
      ic_tag_valid_out_0_51 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6370) begin
      ic_tag_valid_out_0_52 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6385) begin
      ic_tag_valid_out_0_53 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6400) begin
      ic_tag_valid_out_0_54 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6415) begin
      ic_tag_valid_out_0_55 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6430) begin
      ic_tag_valid_out_0_56 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6445) begin
      ic_tag_valid_out_0_57 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6460) begin
      ic_tag_valid_out_0_58 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6475) begin
      ic_tag_valid_out_0_59 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6490) begin
      ic_tag_valid_out_0_60 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6505) begin
      ic_tag_valid_out_0_61 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6520) begin
      ic_tag_valid_out_0_62 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6535) begin
      ic_tag_valid_out_0_63 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7030) begin
      ic_tag_valid_out_0_64 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7045) begin
      ic_tag_valid_out_0_65 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7060) begin
      ic_tag_valid_out_0_66 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7075) begin
      ic_tag_valid_out_0_67 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7090) begin
      ic_tag_valid_out_0_68 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7105) begin
      ic_tag_valid_out_0_69 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7120) begin
      ic_tag_valid_out_0_70 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7135) begin
      ic_tag_valid_out_0_71 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7150) begin
      ic_tag_valid_out_0_72 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7165) begin
      ic_tag_valid_out_0_73 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7180) begin
      ic_tag_valid_out_0_74 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7195) begin
      ic_tag_valid_out_0_75 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7210) begin
      ic_tag_valid_out_0_76 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7225) begin
      ic_tag_valid_out_0_77 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7240) begin
      ic_tag_valid_out_0_78 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7255) begin
      ic_tag_valid_out_0_79 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7270) begin
      ic_tag_valid_out_0_80 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7285) begin
      ic_tag_valid_out_0_81 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7300) begin
      ic_tag_valid_out_0_82 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7315) begin
      ic_tag_valid_out_0_83 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7330) begin
      ic_tag_valid_out_0_84 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7345) begin
      ic_tag_valid_out_0_85 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7360) begin
      ic_tag_valid_out_0_86 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7375) begin
      ic_tag_valid_out_0_87 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7390) begin
      ic_tag_valid_out_0_88 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7405) begin
      ic_tag_valid_out_0_89 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7420) begin
      ic_tag_valid_out_0_90 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7435) begin
      ic_tag_valid_out_0_91 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7450) begin
      ic_tag_valid_out_0_92 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7465) begin
      ic_tag_valid_out_0_93 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7480) begin
      ic_tag_valid_out_0_94 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7495) begin
      ic_tag_valid_out_0_95 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_7990) begin
      ic_tag_valid_out_0_96 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8005) begin
      ic_tag_valid_out_0_97 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8020) begin
      ic_tag_valid_out_0_98 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8035) begin
      ic_tag_valid_out_0_99 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8050) begin
      ic_tag_valid_out_0_100 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8065) begin
      ic_tag_valid_out_0_101 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8080) begin
      ic_tag_valid_out_0_102 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8095) begin
      ic_tag_valid_out_0_103 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8110) begin
      ic_tag_valid_out_0_104 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8125) begin
      ic_tag_valid_out_0_105 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8140) begin
      ic_tag_valid_out_0_106 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8155) begin
      ic_tag_valid_out_0_107 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8170) begin
      ic_tag_valid_out_0_108 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8185) begin
      ic_tag_valid_out_0_109 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8200) begin
      ic_tag_valid_out_0_110 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8215) begin
      ic_tag_valid_out_0_111 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8230) begin
      ic_tag_valid_out_0_112 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8245) begin
      ic_tag_valid_out_0_113 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8260) begin
      ic_tag_valid_out_0_114 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8275) begin
      ic_tag_valid_out_0_115 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8290) begin
      ic_tag_valid_out_0_116 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8305) begin
      ic_tag_valid_out_0_117 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8320) begin
      ic_tag_valid_out_0_118 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8335) begin
      ic_tag_valid_out_0_119 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8350) begin
      ic_tag_valid_out_0_120 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8365) begin
      ic_tag_valid_out_0_121 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8380) begin
      ic_tag_valid_out_0_122 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8395) begin
      ic_tag_valid_out_0_123 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8410) begin
      ic_tag_valid_out_0_124 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8425) begin
      ic_tag_valid_out_0_125 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8440) begin
      ic_tag_valid_out_0_126 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8455) begin
      ic_tag_valid_out_0_127 <= _T_5102;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_1211 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1211 <= _T_1210;
    end else begin
      _T_1211 <= io_ic_debug_rd_data;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_memory_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_memory_f <= _T_9834 & io_ifc_fetch_req_bf;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      perr_ic_index_ff <= 7'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= perr_state == 3'h4;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_cmd_req_hold <= 1'h0;
    end else begin
      bus_cmd_req_hold <= _T_2554 & _T_2573;
    end
  end
  always @(posedge rvclkhdr_69_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else begin
      ifu_bus_cmd_valid <= _T_2544 & _T_2550;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (bus_cmd_beat_en) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= _T_2649 & _T_2650;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3880;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rtag_temp <= 3'h0;
    end else begin
      iccm_dma_rtag_temp <= dma_mem_tag_ff;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_temp <= 1'h0;
    end else begin
      iccm_dma_rvalid_temp <= iccm_dma_rvalid_in;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_ecc_error <= 1'h0;
    end else begin
      iccm_dma_ecc_error <= |iccm_double_ecc_error;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rdata_temp <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata_temp <= _T_3054;
    end else begin
      iccm_dma_rdata_temp <= _T_3055;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3876;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= _T_3871 & _T_319;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3945) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en | _T_3948;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      way_status_new_ff <= 1'h0;
    end else if (_T_3948) begin
      way_status_new_ff <= io_ic_debug_wr_data[4];
    end else if (_T_9725) begin
      way_status_new_ff <= replace_way_mb_any_0;
    end else begin
      way_status_new_ff <= way_status_hit_new;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren | ic_debug_tag_wr_en;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3948) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9747 <= 1'h0;
    end else begin
      _T_9747 <= _T_233 & _T_209;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9748 <= 1'h0;
    end else begin
      _T_9748 <= _T_225 & _T_247;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9749 <= 1'h0;
    end else begin
      _T_9749 <= ic_byp_hit_f & ifu_byp_data_err_new;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9753 <= 1'h0;
    end else begin
      _T_9753 <= _T_9751 & miss_pending;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9754 <= 1'h0;
    end else begin
      _T_9754 <= _T_2568 & _T_2573;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_9775 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_9775 <= ic_debug_rd_en_ff;
    end
  end
endmodule
