module el2_dec_trigger(
  input         clock,
  input         reset,
  input         io_trigger_pkt_any_0_select,
  input         io_trigger_pkt_any_0_match_,
  input         io_trigger_pkt_any_0_store,
  input         io_trigger_pkt_any_0_load,
  input         io_trigger_pkt_any_0_execute,
  input         io_trigger_pkt_any_0_m,
  input  [31:0] io_trigger_pkt_any_0_tdata2,
  input         io_trigger_pkt_any_1_select,
  input         io_trigger_pkt_any_1_match_,
  input         io_trigger_pkt_any_1_store,
  input         io_trigger_pkt_any_1_load,
  input         io_trigger_pkt_any_1_execute,
  input         io_trigger_pkt_any_1_m,
  input  [31:0] io_trigger_pkt_any_1_tdata2,
  input         io_trigger_pkt_any_2_select,
  input         io_trigger_pkt_any_2_match_,
  input         io_trigger_pkt_any_2_store,
  input         io_trigger_pkt_any_2_load,
  input         io_trigger_pkt_any_2_execute,
  input         io_trigger_pkt_any_2_m,
  input  [31:0] io_trigger_pkt_any_2_tdata2,
  input         io_trigger_pkt_any_3_select,
  input         io_trigger_pkt_any_3_match_,
  input         io_trigger_pkt_any_3_store,
  input         io_trigger_pkt_any_3_load,
  input         io_trigger_pkt_any_3_execute,
  input         io_trigger_pkt_any_3_m,
  input  [31:0] io_trigger_pkt_any_3_tdata2,
  input  [30:0] io_dec_i0_pc_d,
  output [3:0]  io_dec_i0_trigger_match_d
);
  wire  _T = ~io_trigger_pkt_any_0_select; // @[el2_dec_trigger.scala 14:63]
  wire  _T_1 = _T & io_trigger_pkt_any_0_execute; // @[el2_dec_trigger.scala 14:93]
  wire [9:0] _T_11 = {_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [18:0] _T_20 = {_T_11,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [27:0] _T_29 = {_T_20,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [31:0] _T_33 = {_T_29,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [31:0] _T_35 = {io_dec_i0_pc_d,io_trigger_pkt_any_0_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_0 = _T_33 & _T_35; // @[el2_dec_trigger.scala 14:127]
  wire  _T_37 = ~io_trigger_pkt_any_1_select; // @[el2_dec_trigger.scala 14:63]
  wire  _T_38 = _T_37 & io_trigger_pkt_any_1_execute; // @[el2_dec_trigger.scala 14:93]
  wire [9:0] _T_48 = {_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [18:0] _T_57 = {_T_48,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [27:0] _T_66 = {_T_57,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [31:0] _T_70 = {_T_66,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [31:0] _T_72 = {io_dec_i0_pc_d,io_trigger_pkt_any_1_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_1 = _T_70 & _T_72; // @[el2_dec_trigger.scala 14:127]
  wire  _T_74 = ~io_trigger_pkt_any_2_select; // @[el2_dec_trigger.scala 14:63]
  wire  _T_75 = _T_74 & io_trigger_pkt_any_2_execute; // @[el2_dec_trigger.scala 14:93]
  wire [9:0] _T_85 = {_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [18:0] _T_94 = {_T_85,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [27:0] _T_103 = {_T_94,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [31:0] _T_107 = {_T_103,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [31:0] _T_109 = {io_dec_i0_pc_d,io_trigger_pkt_any_2_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_2 = _T_107 & _T_109; // @[el2_dec_trigger.scala 14:127]
  wire  _T_111 = ~io_trigger_pkt_any_3_select; // @[el2_dec_trigger.scala 14:63]
  wire  _T_112 = _T_111 & io_trigger_pkt_any_3_execute; // @[el2_dec_trigger.scala 14:93]
  wire [9:0] _T_122 = {_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [18:0] _T_131 = {_T_122,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [27:0] _T_140 = {_T_131,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [31:0] _T_144 = {_T_140,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [31:0] _T_146 = {io_dec_i0_pc_d,io_trigger_pkt_any_3_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_3 = _T_144 & _T_146; // @[el2_dec_trigger.scala 14:127]
  wire  _T_148 = io_trigger_pkt_any_0_execute & io_trigger_pkt_any_0_m; // @[el2_dec_trigger.scala 15:83]
  wire  _T_153 = &io_trigger_pkt_any_0_tdata2; // @[el2_lib.scala 216:73]
  wire  _T_154 = ~_T_153; // @[el2_lib.scala 216:47]
  wire  _T_155 = io_trigger_pkt_any_0_match_ & _T_154; // @[el2_lib.scala 216:44]
  wire  _T_158 = io_trigger_pkt_any_0_tdata2[0] == dec_i0_match_data_0[0]; // @[el2_lib.scala 217:52]
  wire  _T_159 = _T_155 | _T_158; // @[el2_lib.scala 217:41]
  wire  _T_161 = &io_trigger_pkt_any_0_tdata2[0]; // @[el2_lib.scala 219:37]
  wire  _T_162 = _T_161 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_165 = io_trigger_pkt_any_0_tdata2[1] == dec_i0_match_data_0[1]; // @[el2_lib.scala 219:79]
  wire  _T_166 = _T_162 | _T_165; // @[el2_lib.scala 219:24]
  wire  _T_168 = &io_trigger_pkt_any_0_tdata2[1:0]; // @[el2_lib.scala 219:37]
  wire  _T_169 = _T_168 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_172 = io_trigger_pkt_any_0_tdata2[2] == dec_i0_match_data_0[2]; // @[el2_lib.scala 219:79]
  wire  _T_173 = _T_169 | _T_172; // @[el2_lib.scala 219:24]
  wire  _T_175 = &io_trigger_pkt_any_0_tdata2[2:0]; // @[el2_lib.scala 219:37]
  wire  _T_176 = _T_175 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_179 = io_trigger_pkt_any_0_tdata2[3] == dec_i0_match_data_0[3]; // @[el2_lib.scala 219:79]
  wire  _T_180 = _T_176 | _T_179; // @[el2_lib.scala 219:24]
  wire  _T_182 = &io_trigger_pkt_any_0_tdata2[3:0]; // @[el2_lib.scala 219:37]
  wire  _T_183 = _T_182 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_186 = io_trigger_pkt_any_0_tdata2[4] == dec_i0_match_data_0[4]; // @[el2_lib.scala 219:79]
  wire  _T_187 = _T_183 | _T_186; // @[el2_lib.scala 219:24]
  wire  _T_189 = &io_trigger_pkt_any_0_tdata2[4:0]; // @[el2_lib.scala 219:37]
  wire  _T_190 = _T_189 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_193 = io_trigger_pkt_any_0_tdata2[5] == dec_i0_match_data_0[5]; // @[el2_lib.scala 219:79]
  wire  _T_194 = _T_190 | _T_193; // @[el2_lib.scala 219:24]
  wire  _T_196 = &io_trigger_pkt_any_0_tdata2[5:0]; // @[el2_lib.scala 219:37]
  wire  _T_197 = _T_196 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_200 = io_trigger_pkt_any_0_tdata2[6] == dec_i0_match_data_0[6]; // @[el2_lib.scala 219:79]
  wire  _T_201 = _T_197 | _T_200; // @[el2_lib.scala 219:24]
  wire  _T_203 = &io_trigger_pkt_any_0_tdata2[6:0]; // @[el2_lib.scala 219:37]
  wire  _T_204 = _T_203 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_207 = io_trigger_pkt_any_0_tdata2[7] == dec_i0_match_data_0[7]; // @[el2_lib.scala 219:79]
  wire  _T_208 = _T_204 | _T_207; // @[el2_lib.scala 219:24]
  wire  _T_210 = &io_trigger_pkt_any_0_tdata2[7:0]; // @[el2_lib.scala 219:37]
  wire  _T_211 = _T_210 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_214 = io_trigger_pkt_any_0_tdata2[8] == dec_i0_match_data_0[8]; // @[el2_lib.scala 219:79]
  wire  _T_215 = _T_211 | _T_214; // @[el2_lib.scala 219:24]
  wire  _T_217 = &io_trigger_pkt_any_0_tdata2[8:0]; // @[el2_lib.scala 219:37]
  wire  _T_218 = _T_217 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_221 = io_trigger_pkt_any_0_tdata2[9] == dec_i0_match_data_0[9]; // @[el2_lib.scala 219:79]
  wire  _T_222 = _T_218 | _T_221; // @[el2_lib.scala 219:24]
  wire  _T_224 = &io_trigger_pkt_any_0_tdata2[9:0]; // @[el2_lib.scala 219:37]
  wire  _T_225 = _T_224 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_228 = io_trigger_pkt_any_0_tdata2[10] == dec_i0_match_data_0[10]; // @[el2_lib.scala 219:79]
  wire  _T_229 = _T_225 | _T_228; // @[el2_lib.scala 219:24]
  wire  _T_231 = &io_trigger_pkt_any_0_tdata2[10:0]; // @[el2_lib.scala 219:37]
  wire  _T_232 = _T_231 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_235 = io_trigger_pkt_any_0_tdata2[11] == dec_i0_match_data_0[11]; // @[el2_lib.scala 219:79]
  wire  _T_236 = _T_232 | _T_235; // @[el2_lib.scala 219:24]
  wire  _T_238 = &io_trigger_pkt_any_0_tdata2[11:0]; // @[el2_lib.scala 219:37]
  wire  _T_239 = _T_238 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_242 = io_trigger_pkt_any_0_tdata2[12] == dec_i0_match_data_0[12]; // @[el2_lib.scala 219:79]
  wire  _T_243 = _T_239 | _T_242; // @[el2_lib.scala 219:24]
  wire  _T_245 = &io_trigger_pkt_any_0_tdata2[12:0]; // @[el2_lib.scala 219:37]
  wire  _T_246 = _T_245 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_249 = io_trigger_pkt_any_0_tdata2[13] == dec_i0_match_data_0[13]; // @[el2_lib.scala 219:79]
  wire  _T_250 = _T_246 | _T_249; // @[el2_lib.scala 219:24]
  wire  _T_252 = &io_trigger_pkt_any_0_tdata2[13:0]; // @[el2_lib.scala 219:37]
  wire  _T_253 = _T_252 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_256 = io_trigger_pkt_any_0_tdata2[14] == dec_i0_match_data_0[14]; // @[el2_lib.scala 219:79]
  wire  _T_257 = _T_253 | _T_256; // @[el2_lib.scala 219:24]
  wire  _T_259 = &io_trigger_pkt_any_0_tdata2[14:0]; // @[el2_lib.scala 219:37]
  wire  _T_260 = _T_259 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_263 = io_trigger_pkt_any_0_tdata2[15] == dec_i0_match_data_0[15]; // @[el2_lib.scala 219:79]
  wire  _T_264 = _T_260 | _T_263; // @[el2_lib.scala 219:24]
  wire  _T_266 = &io_trigger_pkt_any_0_tdata2[15:0]; // @[el2_lib.scala 219:37]
  wire  _T_267 = _T_266 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_270 = io_trigger_pkt_any_0_tdata2[16] == dec_i0_match_data_0[16]; // @[el2_lib.scala 219:79]
  wire  _T_271 = _T_267 | _T_270; // @[el2_lib.scala 219:24]
  wire  _T_273 = &io_trigger_pkt_any_0_tdata2[16:0]; // @[el2_lib.scala 219:37]
  wire  _T_274 = _T_273 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_277 = io_trigger_pkt_any_0_tdata2[17] == dec_i0_match_data_0[17]; // @[el2_lib.scala 219:79]
  wire  _T_278 = _T_274 | _T_277; // @[el2_lib.scala 219:24]
  wire  _T_280 = &io_trigger_pkt_any_0_tdata2[17:0]; // @[el2_lib.scala 219:37]
  wire  _T_281 = _T_280 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_284 = io_trigger_pkt_any_0_tdata2[18] == dec_i0_match_data_0[18]; // @[el2_lib.scala 219:79]
  wire  _T_285 = _T_281 | _T_284; // @[el2_lib.scala 219:24]
  wire  _T_287 = &io_trigger_pkt_any_0_tdata2[18:0]; // @[el2_lib.scala 219:37]
  wire  _T_288 = _T_287 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_291 = io_trigger_pkt_any_0_tdata2[19] == dec_i0_match_data_0[19]; // @[el2_lib.scala 219:79]
  wire  _T_292 = _T_288 | _T_291; // @[el2_lib.scala 219:24]
  wire  _T_294 = &io_trigger_pkt_any_0_tdata2[19:0]; // @[el2_lib.scala 219:37]
  wire  _T_295 = _T_294 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_298 = io_trigger_pkt_any_0_tdata2[20] == dec_i0_match_data_0[20]; // @[el2_lib.scala 219:79]
  wire  _T_299 = _T_295 | _T_298; // @[el2_lib.scala 219:24]
  wire  _T_301 = &io_trigger_pkt_any_0_tdata2[20:0]; // @[el2_lib.scala 219:37]
  wire  _T_302 = _T_301 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_305 = io_trigger_pkt_any_0_tdata2[21] == dec_i0_match_data_0[21]; // @[el2_lib.scala 219:79]
  wire  _T_306 = _T_302 | _T_305; // @[el2_lib.scala 219:24]
  wire  _T_308 = &io_trigger_pkt_any_0_tdata2[21:0]; // @[el2_lib.scala 219:37]
  wire  _T_309 = _T_308 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_312 = io_trigger_pkt_any_0_tdata2[22] == dec_i0_match_data_0[22]; // @[el2_lib.scala 219:79]
  wire  _T_313 = _T_309 | _T_312; // @[el2_lib.scala 219:24]
  wire  _T_315 = &io_trigger_pkt_any_0_tdata2[22:0]; // @[el2_lib.scala 219:37]
  wire  _T_316 = _T_315 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_319 = io_trigger_pkt_any_0_tdata2[23] == dec_i0_match_data_0[23]; // @[el2_lib.scala 219:79]
  wire  _T_320 = _T_316 | _T_319; // @[el2_lib.scala 219:24]
  wire  _T_322 = &io_trigger_pkt_any_0_tdata2[23:0]; // @[el2_lib.scala 219:37]
  wire  _T_323 = _T_322 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_326 = io_trigger_pkt_any_0_tdata2[24] == dec_i0_match_data_0[24]; // @[el2_lib.scala 219:79]
  wire  _T_327 = _T_323 | _T_326; // @[el2_lib.scala 219:24]
  wire  _T_329 = &io_trigger_pkt_any_0_tdata2[24:0]; // @[el2_lib.scala 219:37]
  wire  _T_330 = _T_329 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_333 = io_trigger_pkt_any_0_tdata2[25] == dec_i0_match_data_0[25]; // @[el2_lib.scala 219:79]
  wire  _T_334 = _T_330 | _T_333; // @[el2_lib.scala 219:24]
  wire  _T_336 = &io_trigger_pkt_any_0_tdata2[25:0]; // @[el2_lib.scala 219:37]
  wire  _T_337 = _T_336 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_340 = io_trigger_pkt_any_0_tdata2[26] == dec_i0_match_data_0[26]; // @[el2_lib.scala 219:79]
  wire  _T_341 = _T_337 | _T_340; // @[el2_lib.scala 219:24]
  wire  _T_343 = &io_trigger_pkt_any_0_tdata2[26:0]; // @[el2_lib.scala 219:37]
  wire  _T_344 = _T_343 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_347 = io_trigger_pkt_any_0_tdata2[27] == dec_i0_match_data_0[27]; // @[el2_lib.scala 219:79]
  wire  _T_348 = _T_344 | _T_347; // @[el2_lib.scala 219:24]
  wire  _T_350 = &io_trigger_pkt_any_0_tdata2[27:0]; // @[el2_lib.scala 219:37]
  wire  _T_351 = _T_350 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_354 = io_trigger_pkt_any_0_tdata2[28] == dec_i0_match_data_0[28]; // @[el2_lib.scala 219:79]
  wire  _T_355 = _T_351 | _T_354; // @[el2_lib.scala 219:24]
  wire  _T_357 = &io_trigger_pkt_any_0_tdata2[28:0]; // @[el2_lib.scala 219:37]
  wire  _T_358 = _T_357 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_361 = io_trigger_pkt_any_0_tdata2[29] == dec_i0_match_data_0[29]; // @[el2_lib.scala 219:79]
  wire  _T_362 = _T_358 | _T_361; // @[el2_lib.scala 219:24]
  wire  _T_364 = &io_trigger_pkt_any_0_tdata2[29:0]; // @[el2_lib.scala 219:37]
  wire  _T_365 = _T_364 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_368 = io_trigger_pkt_any_0_tdata2[30] == dec_i0_match_data_0[30]; // @[el2_lib.scala 219:79]
  wire  _T_369 = _T_365 | _T_368; // @[el2_lib.scala 219:24]
  wire  _T_371 = &io_trigger_pkt_any_0_tdata2[30:0]; // @[el2_lib.scala 219:37]
  wire  _T_372 = _T_371 & _T_155; // @[el2_lib.scala 219:42]
  wire  _T_375 = io_trigger_pkt_any_0_tdata2[31] == dec_i0_match_data_0[31]; // @[el2_lib.scala 219:79]
  wire  _T_376 = _T_372 | _T_375; // @[el2_lib.scala 219:24]
  wire [7:0] _T_383 = {_T_208,_T_201,_T_194,_T_187,_T_180,_T_173,_T_166,_T_159}; // @[el2_lib.scala 220:14]
  wire [15:0] _T_391 = {_T_264,_T_257,_T_250,_T_243,_T_236,_T_229,_T_222,_T_215,_T_383}; // @[el2_lib.scala 220:14]
  wire [7:0] _T_398 = {_T_320,_T_313,_T_306,_T_299,_T_292,_T_285,_T_278,_T_271}; // @[el2_lib.scala 220:14]
  wire [31:0] _T_407 = {_T_376,_T_369,_T_362,_T_355,_T_348,_T_341,_T_334,_T_327,_T_398,_T_391}; // @[el2_lib.scala 220:14]
  wire  _T_408 = &_T_407; // @[el2_lib.scala 220:21]
  wire  _T_409 = _T_148 & _T_408; // @[el2_dec_trigger.scala 15:109]
  wire  _T_410 = io_trigger_pkt_any_1_execute & io_trigger_pkt_any_1_m; // @[el2_dec_trigger.scala 15:83]
  wire  _T_415 = &io_trigger_pkt_any_1_tdata2; // @[el2_lib.scala 216:73]
  wire  _T_416 = ~_T_415; // @[el2_lib.scala 216:47]
  wire  _T_417 = io_trigger_pkt_any_1_match_ & _T_416; // @[el2_lib.scala 216:44]
  wire  _T_420 = io_trigger_pkt_any_1_tdata2[0] == dec_i0_match_data_1[0]; // @[el2_lib.scala 217:52]
  wire  _T_421 = _T_417 | _T_420; // @[el2_lib.scala 217:41]
  wire  _T_423 = &io_trigger_pkt_any_1_tdata2[0]; // @[el2_lib.scala 219:37]
  wire  _T_424 = _T_423 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_427 = io_trigger_pkt_any_1_tdata2[1] == dec_i0_match_data_1[1]; // @[el2_lib.scala 219:79]
  wire  _T_428 = _T_424 | _T_427; // @[el2_lib.scala 219:24]
  wire  _T_430 = &io_trigger_pkt_any_1_tdata2[1:0]; // @[el2_lib.scala 219:37]
  wire  _T_431 = _T_430 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_434 = io_trigger_pkt_any_1_tdata2[2] == dec_i0_match_data_1[2]; // @[el2_lib.scala 219:79]
  wire  _T_435 = _T_431 | _T_434; // @[el2_lib.scala 219:24]
  wire  _T_437 = &io_trigger_pkt_any_1_tdata2[2:0]; // @[el2_lib.scala 219:37]
  wire  _T_438 = _T_437 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_441 = io_trigger_pkt_any_1_tdata2[3] == dec_i0_match_data_1[3]; // @[el2_lib.scala 219:79]
  wire  _T_442 = _T_438 | _T_441; // @[el2_lib.scala 219:24]
  wire  _T_444 = &io_trigger_pkt_any_1_tdata2[3:0]; // @[el2_lib.scala 219:37]
  wire  _T_445 = _T_444 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_448 = io_trigger_pkt_any_1_tdata2[4] == dec_i0_match_data_1[4]; // @[el2_lib.scala 219:79]
  wire  _T_449 = _T_445 | _T_448; // @[el2_lib.scala 219:24]
  wire  _T_451 = &io_trigger_pkt_any_1_tdata2[4:0]; // @[el2_lib.scala 219:37]
  wire  _T_452 = _T_451 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_455 = io_trigger_pkt_any_1_tdata2[5] == dec_i0_match_data_1[5]; // @[el2_lib.scala 219:79]
  wire  _T_456 = _T_452 | _T_455; // @[el2_lib.scala 219:24]
  wire  _T_458 = &io_trigger_pkt_any_1_tdata2[5:0]; // @[el2_lib.scala 219:37]
  wire  _T_459 = _T_458 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_462 = io_trigger_pkt_any_1_tdata2[6] == dec_i0_match_data_1[6]; // @[el2_lib.scala 219:79]
  wire  _T_463 = _T_459 | _T_462; // @[el2_lib.scala 219:24]
  wire  _T_465 = &io_trigger_pkt_any_1_tdata2[6:0]; // @[el2_lib.scala 219:37]
  wire  _T_466 = _T_465 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_469 = io_trigger_pkt_any_1_tdata2[7] == dec_i0_match_data_1[7]; // @[el2_lib.scala 219:79]
  wire  _T_470 = _T_466 | _T_469; // @[el2_lib.scala 219:24]
  wire  _T_472 = &io_trigger_pkt_any_1_tdata2[7:0]; // @[el2_lib.scala 219:37]
  wire  _T_473 = _T_472 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_476 = io_trigger_pkt_any_1_tdata2[8] == dec_i0_match_data_1[8]; // @[el2_lib.scala 219:79]
  wire  _T_477 = _T_473 | _T_476; // @[el2_lib.scala 219:24]
  wire  _T_479 = &io_trigger_pkt_any_1_tdata2[8:0]; // @[el2_lib.scala 219:37]
  wire  _T_480 = _T_479 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_483 = io_trigger_pkt_any_1_tdata2[9] == dec_i0_match_data_1[9]; // @[el2_lib.scala 219:79]
  wire  _T_484 = _T_480 | _T_483; // @[el2_lib.scala 219:24]
  wire  _T_486 = &io_trigger_pkt_any_1_tdata2[9:0]; // @[el2_lib.scala 219:37]
  wire  _T_487 = _T_486 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_490 = io_trigger_pkt_any_1_tdata2[10] == dec_i0_match_data_1[10]; // @[el2_lib.scala 219:79]
  wire  _T_491 = _T_487 | _T_490; // @[el2_lib.scala 219:24]
  wire  _T_493 = &io_trigger_pkt_any_1_tdata2[10:0]; // @[el2_lib.scala 219:37]
  wire  _T_494 = _T_493 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_497 = io_trigger_pkt_any_1_tdata2[11] == dec_i0_match_data_1[11]; // @[el2_lib.scala 219:79]
  wire  _T_498 = _T_494 | _T_497; // @[el2_lib.scala 219:24]
  wire  _T_500 = &io_trigger_pkt_any_1_tdata2[11:0]; // @[el2_lib.scala 219:37]
  wire  _T_501 = _T_500 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_504 = io_trigger_pkt_any_1_tdata2[12] == dec_i0_match_data_1[12]; // @[el2_lib.scala 219:79]
  wire  _T_505 = _T_501 | _T_504; // @[el2_lib.scala 219:24]
  wire  _T_507 = &io_trigger_pkt_any_1_tdata2[12:0]; // @[el2_lib.scala 219:37]
  wire  _T_508 = _T_507 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_511 = io_trigger_pkt_any_1_tdata2[13] == dec_i0_match_data_1[13]; // @[el2_lib.scala 219:79]
  wire  _T_512 = _T_508 | _T_511; // @[el2_lib.scala 219:24]
  wire  _T_514 = &io_trigger_pkt_any_1_tdata2[13:0]; // @[el2_lib.scala 219:37]
  wire  _T_515 = _T_514 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_518 = io_trigger_pkt_any_1_tdata2[14] == dec_i0_match_data_1[14]; // @[el2_lib.scala 219:79]
  wire  _T_519 = _T_515 | _T_518; // @[el2_lib.scala 219:24]
  wire  _T_521 = &io_trigger_pkt_any_1_tdata2[14:0]; // @[el2_lib.scala 219:37]
  wire  _T_522 = _T_521 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_525 = io_trigger_pkt_any_1_tdata2[15] == dec_i0_match_data_1[15]; // @[el2_lib.scala 219:79]
  wire  _T_526 = _T_522 | _T_525; // @[el2_lib.scala 219:24]
  wire  _T_528 = &io_trigger_pkt_any_1_tdata2[15:0]; // @[el2_lib.scala 219:37]
  wire  _T_529 = _T_528 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_532 = io_trigger_pkt_any_1_tdata2[16] == dec_i0_match_data_1[16]; // @[el2_lib.scala 219:79]
  wire  _T_533 = _T_529 | _T_532; // @[el2_lib.scala 219:24]
  wire  _T_535 = &io_trigger_pkt_any_1_tdata2[16:0]; // @[el2_lib.scala 219:37]
  wire  _T_536 = _T_535 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_539 = io_trigger_pkt_any_1_tdata2[17] == dec_i0_match_data_1[17]; // @[el2_lib.scala 219:79]
  wire  _T_540 = _T_536 | _T_539; // @[el2_lib.scala 219:24]
  wire  _T_542 = &io_trigger_pkt_any_1_tdata2[17:0]; // @[el2_lib.scala 219:37]
  wire  _T_543 = _T_542 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_546 = io_trigger_pkt_any_1_tdata2[18] == dec_i0_match_data_1[18]; // @[el2_lib.scala 219:79]
  wire  _T_547 = _T_543 | _T_546; // @[el2_lib.scala 219:24]
  wire  _T_549 = &io_trigger_pkt_any_1_tdata2[18:0]; // @[el2_lib.scala 219:37]
  wire  _T_550 = _T_549 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_553 = io_trigger_pkt_any_1_tdata2[19] == dec_i0_match_data_1[19]; // @[el2_lib.scala 219:79]
  wire  _T_554 = _T_550 | _T_553; // @[el2_lib.scala 219:24]
  wire  _T_556 = &io_trigger_pkt_any_1_tdata2[19:0]; // @[el2_lib.scala 219:37]
  wire  _T_557 = _T_556 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_560 = io_trigger_pkt_any_1_tdata2[20] == dec_i0_match_data_1[20]; // @[el2_lib.scala 219:79]
  wire  _T_561 = _T_557 | _T_560; // @[el2_lib.scala 219:24]
  wire  _T_563 = &io_trigger_pkt_any_1_tdata2[20:0]; // @[el2_lib.scala 219:37]
  wire  _T_564 = _T_563 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_567 = io_trigger_pkt_any_1_tdata2[21] == dec_i0_match_data_1[21]; // @[el2_lib.scala 219:79]
  wire  _T_568 = _T_564 | _T_567; // @[el2_lib.scala 219:24]
  wire  _T_570 = &io_trigger_pkt_any_1_tdata2[21:0]; // @[el2_lib.scala 219:37]
  wire  _T_571 = _T_570 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_574 = io_trigger_pkt_any_1_tdata2[22] == dec_i0_match_data_1[22]; // @[el2_lib.scala 219:79]
  wire  _T_575 = _T_571 | _T_574; // @[el2_lib.scala 219:24]
  wire  _T_577 = &io_trigger_pkt_any_1_tdata2[22:0]; // @[el2_lib.scala 219:37]
  wire  _T_578 = _T_577 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_581 = io_trigger_pkt_any_1_tdata2[23] == dec_i0_match_data_1[23]; // @[el2_lib.scala 219:79]
  wire  _T_582 = _T_578 | _T_581; // @[el2_lib.scala 219:24]
  wire  _T_584 = &io_trigger_pkt_any_1_tdata2[23:0]; // @[el2_lib.scala 219:37]
  wire  _T_585 = _T_584 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_588 = io_trigger_pkt_any_1_tdata2[24] == dec_i0_match_data_1[24]; // @[el2_lib.scala 219:79]
  wire  _T_589 = _T_585 | _T_588; // @[el2_lib.scala 219:24]
  wire  _T_591 = &io_trigger_pkt_any_1_tdata2[24:0]; // @[el2_lib.scala 219:37]
  wire  _T_592 = _T_591 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_595 = io_trigger_pkt_any_1_tdata2[25] == dec_i0_match_data_1[25]; // @[el2_lib.scala 219:79]
  wire  _T_596 = _T_592 | _T_595; // @[el2_lib.scala 219:24]
  wire  _T_598 = &io_trigger_pkt_any_1_tdata2[25:0]; // @[el2_lib.scala 219:37]
  wire  _T_599 = _T_598 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_602 = io_trigger_pkt_any_1_tdata2[26] == dec_i0_match_data_1[26]; // @[el2_lib.scala 219:79]
  wire  _T_603 = _T_599 | _T_602; // @[el2_lib.scala 219:24]
  wire  _T_605 = &io_trigger_pkt_any_1_tdata2[26:0]; // @[el2_lib.scala 219:37]
  wire  _T_606 = _T_605 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_609 = io_trigger_pkt_any_1_tdata2[27] == dec_i0_match_data_1[27]; // @[el2_lib.scala 219:79]
  wire  _T_610 = _T_606 | _T_609; // @[el2_lib.scala 219:24]
  wire  _T_612 = &io_trigger_pkt_any_1_tdata2[27:0]; // @[el2_lib.scala 219:37]
  wire  _T_613 = _T_612 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_616 = io_trigger_pkt_any_1_tdata2[28] == dec_i0_match_data_1[28]; // @[el2_lib.scala 219:79]
  wire  _T_617 = _T_613 | _T_616; // @[el2_lib.scala 219:24]
  wire  _T_619 = &io_trigger_pkt_any_1_tdata2[28:0]; // @[el2_lib.scala 219:37]
  wire  _T_620 = _T_619 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_623 = io_trigger_pkt_any_1_tdata2[29] == dec_i0_match_data_1[29]; // @[el2_lib.scala 219:79]
  wire  _T_624 = _T_620 | _T_623; // @[el2_lib.scala 219:24]
  wire  _T_626 = &io_trigger_pkt_any_1_tdata2[29:0]; // @[el2_lib.scala 219:37]
  wire  _T_627 = _T_626 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_630 = io_trigger_pkt_any_1_tdata2[30] == dec_i0_match_data_1[30]; // @[el2_lib.scala 219:79]
  wire  _T_631 = _T_627 | _T_630; // @[el2_lib.scala 219:24]
  wire  _T_633 = &io_trigger_pkt_any_1_tdata2[30:0]; // @[el2_lib.scala 219:37]
  wire  _T_634 = _T_633 & _T_417; // @[el2_lib.scala 219:42]
  wire  _T_637 = io_trigger_pkt_any_1_tdata2[31] == dec_i0_match_data_1[31]; // @[el2_lib.scala 219:79]
  wire  _T_638 = _T_634 | _T_637; // @[el2_lib.scala 219:24]
  wire [7:0] _T_645 = {_T_470,_T_463,_T_456,_T_449,_T_442,_T_435,_T_428,_T_421}; // @[el2_lib.scala 220:14]
  wire [15:0] _T_653 = {_T_526,_T_519,_T_512,_T_505,_T_498,_T_491,_T_484,_T_477,_T_645}; // @[el2_lib.scala 220:14]
  wire [7:0] _T_660 = {_T_582,_T_575,_T_568,_T_561,_T_554,_T_547,_T_540,_T_533}; // @[el2_lib.scala 220:14]
  wire [31:0] _T_669 = {_T_638,_T_631,_T_624,_T_617,_T_610,_T_603,_T_596,_T_589,_T_660,_T_653}; // @[el2_lib.scala 220:14]
  wire  _T_670 = &_T_669; // @[el2_lib.scala 220:21]
  wire  _T_671 = _T_410 & _T_670; // @[el2_dec_trigger.scala 15:109]
  wire  _T_672 = io_trigger_pkt_any_2_execute & io_trigger_pkt_any_2_m; // @[el2_dec_trigger.scala 15:83]
  wire  _T_677 = &io_trigger_pkt_any_2_tdata2; // @[el2_lib.scala 216:73]
  wire  _T_678 = ~_T_677; // @[el2_lib.scala 216:47]
  wire  _T_679 = io_trigger_pkt_any_2_match_ & _T_678; // @[el2_lib.scala 216:44]
  wire  _T_682 = io_trigger_pkt_any_2_tdata2[0] == dec_i0_match_data_2[0]; // @[el2_lib.scala 217:52]
  wire  _T_683 = _T_679 | _T_682; // @[el2_lib.scala 217:41]
  wire  _T_685 = &io_trigger_pkt_any_2_tdata2[0]; // @[el2_lib.scala 219:37]
  wire  _T_686 = _T_685 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_689 = io_trigger_pkt_any_2_tdata2[1] == dec_i0_match_data_2[1]; // @[el2_lib.scala 219:79]
  wire  _T_690 = _T_686 | _T_689; // @[el2_lib.scala 219:24]
  wire  _T_692 = &io_trigger_pkt_any_2_tdata2[1:0]; // @[el2_lib.scala 219:37]
  wire  _T_693 = _T_692 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_696 = io_trigger_pkt_any_2_tdata2[2] == dec_i0_match_data_2[2]; // @[el2_lib.scala 219:79]
  wire  _T_697 = _T_693 | _T_696; // @[el2_lib.scala 219:24]
  wire  _T_699 = &io_trigger_pkt_any_2_tdata2[2:0]; // @[el2_lib.scala 219:37]
  wire  _T_700 = _T_699 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_703 = io_trigger_pkt_any_2_tdata2[3] == dec_i0_match_data_2[3]; // @[el2_lib.scala 219:79]
  wire  _T_704 = _T_700 | _T_703; // @[el2_lib.scala 219:24]
  wire  _T_706 = &io_trigger_pkt_any_2_tdata2[3:0]; // @[el2_lib.scala 219:37]
  wire  _T_707 = _T_706 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_710 = io_trigger_pkt_any_2_tdata2[4] == dec_i0_match_data_2[4]; // @[el2_lib.scala 219:79]
  wire  _T_711 = _T_707 | _T_710; // @[el2_lib.scala 219:24]
  wire  _T_713 = &io_trigger_pkt_any_2_tdata2[4:0]; // @[el2_lib.scala 219:37]
  wire  _T_714 = _T_713 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_717 = io_trigger_pkt_any_2_tdata2[5] == dec_i0_match_data_2[5]; // @[el2_lib.scala 219:79]
  wire  _T_718 = _T_714 | _T_717; // @[el2_lib.scala 219:24]
  wire  _T_720 = &io_trigger_pkt_any_2_tdata2[5:0]; // @[el2_lib.scala 219:37]
  wire  _T_721 = _T_720 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_724 = io_trigger_pkt_any_2_tdata2[6] == dec_i0_match_data_2[6]; // @[el2_lib.scala 219:79]
  wire  _T_725 = _T_721 | _T_724; // @[el2_lib.scala 219:24]
  wire  _T_727 = &io_trigger_pkt_any_2_tdata2[6:0]; // @[el2_lib.scala 219:37]
  wire  _T_728 = _T_727 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_731 = io_trigger_pkt_any_2_tdata2[7] == dec_i0_match_data_2[7]; // @[el2_lib.scala 219:79]
  wire  _T_732 = _T_728 | _T_731; // @[el2_lib.scala 219:24]
  wire  _T_734 = &io_trigger_pkt_any_2_tdata2[7:0]; // @[el2_lib.scala 219:37]
  wire  _T_735 = _T_734 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_738 = io_trigger_pkt_any_2_tdata2[8] == dec_i0_match_data_2[8]; // @[el2_lib.scala 219:79]
  wire  _T_739 = _T_735 | _T_738; // @[el2_lib.scala 219:24]
  wire  _T_741 = &io_trigger_pkt_any_2_tdata2[8:0]; // @[el2_lib.scala 219:37]
  wire  _T_742 = _T_741 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_745 = io_trigger_pkt_any_2_tdata2[9] == dec_i0_match_data_2[9]; // @[el2_lib.scala 219:79]
  wire  _T_746 = _T_742 | _T_745; // @[el2_lib.scala 219:24]
  wire  _T_748 = &io_trigger_pkt_any_2_tdata2[9:0]; // @[el2_lib.scala 219:37]
  wire  _T_749 = _T_748 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_752 = io_trigger_pkt_any_2_tdata2[10] == dec_i0_match_data_2[10]; // @[el2_lib.scala 219:79]
  wire  _T_753 = _T_749 | _T_752; // @[el2_lib.scala 219:24]
  wire  _T_755 = &io_trigger_pkt_any_2_tdata2[10:0]; // @[el2_lib.scala 219:37]
  wire  _T_756 = _T_755 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_759 = io_trigger_pkt_any_2_tdata2[11] == dec_i0_match_data_2[11]; // @[el2_lib.scala 219:79]
  wire  _T_760 = _T_756 | _T_759; // @[el2_lib.scala 219:24]
  wire  _T_762 = &io_trigger_pkt_any_2_tdata2[11:0]; // @[el2_lib.scala 219:37]
  wire  _T_763 = _T_762 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_766 = io_trigger_pkt_any_2_tdata2[12] == dec_i0_match_data_2[12]; // @[el2_lib.scala 219:79]
  wire  _T_767 = _T_763 | _T_766; // @[el2_lib.scala 219:24]
  wire  _T_769 = &io_trigger_pkt_any_2_tdata2[12:0]; // @[el2_lib.scala 219:37]
  wire  _T_770 = _T_769 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_773 = io_trigger_pkt_any_2_tdata2[13] == dec_i0_match_data_2[13]; // @[el2_lib.scala 219:79]
  wire  _T_774 = _T_770 | _T_773; // @[el2_lib.scala 219:24]
  wire  _T_776 = &io_trigger_pkt_any_2_tdata2[13:0]; // @[el2_lib.scala 219:37]
  wire  _T_777 = _T_776 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_780 = io_trigger_pkt_any_2_tdata2[14] == dec_i0_match_data_2[14]; // @[el2_lib.scala 219:79]
  wire  _T_781 = _T_777 | _T_780; // @[el2_lib.scala 219:24]
  wire  _T_783 = &io_trigger_pkt_any_2_tdata2[14:0]; // @[el2_lib.scala 219:37]
  wire  _T_784 = _T_783 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_787 = io_trigger_pkt_any_2_tdata2[15] == dec_i0_match_data_2[15]; // @[el2_lib.scala 219:79]
  wire  _T_788 = _T_784 | _T_787; // @[el2_lib.scala 219:24]
  wire  _T_790 = &io_trigger_pkt_any_2_tdata2[15:0]; // @[el2_lib.scala 219:37]
  wire  _T_791 = _T_790 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_794 = io_trigger_pkt_any_2_tdata2[16] == dec_i0_match_data_2[16]; // @[el2_lib.scala 219:79]
  wire  _T_795 = _T_791 | _T_794; // @[el2_lib.scala 219:24]
  wire  _T_797 = &io_trigger_pkt_any_2_tdata2[16:0]; // @[el2_lib.scala 219:37]
  wire  _T_798 = _T_797 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_801 = io_trigger_pkt_any_2_tdata2[17] == dec_i0_match_data_2[17]; // @[el2_lib.scala 219:79]
  wire  _T_802 = _T_798 | _T_801; // @[el2_lib.scala 219:24]
  wire  _T_804 = &io_trigger_pkt_any_2_tdata2[17:0]; // @[el2_lib.scala 219:37]
  wire  _T_805 = _T_804 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_808 = io_trigger_pkt_any_2_tdata2[18] == dec_i0_match_data_2[18]; // @[el2_lib.scala 219:79]
  wire  _T_809 = _T_805 | _T_808; // @[el2_lib.scala 219:24]
  wire  _T_811 = &io_trigger_pkt_any_2_tdata2[18:0]; // @[el2_lib.scala 219:37]
  wire  _T_812 = _T_811 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_815 = io_trigger_pkt_any_2_tdata2[19] == dec_i0_match_data_2[19]; // @[el2_lib.scala 219:79]
  wire  _T_816 = _T_812 | _T_815; // @[el2_lib.scala 219:24]
  wire  _T_818 = &io_trigger_pkt_any_2_tdata2[19:0]; // @[el2_lib.scala 219:37]
  wire  _T_819 = _T_818 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_822 = io_trigger_pkt_any_2_tdata2[20] == dec_i0_match_data_2[20]; // @[el2_lib.scala 219:79]
  wire  _T_823 = _T_819 | _T_822; // @[el2_lib.scala 219:24]
  wire  _T_825 = &io_trigger_pkt_any_2_tdata2[20:0]; // @[el2_lib.scala 219:37]
  wire  _T_826 = _T_825 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_829 = io_trigger_pkt_any_2_tdata2[21] == dec_i0_match_data_2[21]; // @[el2_lib.scala 219:79]
  wire  _T_830 = _T_826 | _T_829; // @[el2_lib.scala 219:24]
  wire  _T_832 = &io_trigger_pkt_any_2_tdata2[21:0]; // @[el2_lib.scala 219:37]
  wire  _T_833 = _T_832 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_836 = io_trigger_pkt_any_2_tdata2[22] == dec_i0_match_data_2[22]; // @[el2_lib.scala 219:79]
  wire  _T_837 = _T_833 | _T_836; // @[el2_lib.scala 219:24]
  wire  _T_839 = &io_trigger_pkt_any_2_tdata2[22:0]; // @[el2_lib.scala 219:37]
  wire  _T_840 = _T_839 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_843 = io_trigger_pkt_any_2_tdata2[23] == dec_i0_match_data_2[23]; // @[el2_lib.scala 219:79]
  wire  _T_844 = _T_840 | _T_843; // @[el2_lib.scala 219:24]
  wire  _T_846 = &io_trigger_pkt_any_2_tdata2[23:0]; // @[el2_lib.scala 219:37]
  wire  _T_847 = _T_846 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_850 = io_trigger_pkt_any_2_tdata2[24] == dec_i0_match_data_2[24]; // @[el2_lib.scala 219:79]
  wire  _T_851 = _T_847 | _T_850; // @[el2_lib.scala 219:24]
  wire  _T_853 = &io_trigger_pkt_any_2_tdata2[24:0]; // @[el2_lib.scala 219:37]
  wire  _T_854 = _T_853 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_857 = io_trigger_pkt_any_2_tdata2[25] == dec_i0_match_data_2[25]; // @[el2_lib.scala 219:79]
  wire  _T_858 = _T_854 | _T_857; // @[el2_lib.scala 219:24]
  wire  _T_860 = &io_trigger_pkt_any_2_tdata2[25:0]; // @[el2_lib.scala 219:37]
  wire  _T_861 = _T_860 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_864 = io_trigger_pkt_any_2_tdata2[26] == dec_i0_match_data_2[26]; // @[el2_lib.scala 219:79]
  wire  _T_865 = _T_861 | _T_864; // @[el2_lib.scala 219:24]
  wire  _T_867 = &io_trigger_pkt_any_2_tdata2[26:0]; // @[el2_lib.scala 219:37]
  wire  _T_868 = _T_867 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_871 = io_trigger_pkt_any_2_tdata2[27] == dec_i0_match_data_2[27]; // @[el2_lib.scala 219:79]
  wire  _T_872 = _T_868 | _T_871; // @[el2_lib.scala 219:24]
  wire  _T_874 = &io_trigger_pkt_any_2_tdata2[27:0]; // @[el2_lib.scala 219:37]
  wire  _T_875 = _T_874 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_878 = io_trigger_pkt_any_2_tdata2[28] == dec_i0_match_data_2[28]; // @[el2_lib.scala 219:79]
  wire  _T_879 = _T_875 | _T_878; // @[el2_lib.scala 219:24]
  wire  _T_881 = &io_trigger_pkt_any_2_tdata2[28:0]; // @[el2_lib.scala 219:37]
  wire  _T_882 = _T_881 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_885 = io_trigger_pkt_any_2_tdata2[29] == dec_i0_match_data_2[29]; // @[el2_lib.scala 219:79]
  wire  _T_886 = _T_882 | _T_885; // @[el2_lib.scala 219:24]
  wire  _T_888 = &io_trigger_pkt_any_2_tdata2[29:0]; // @[el2_lib.scala 219:37]
  wire  _T_889 = _T_888 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_892 = io_trigger_pkt_any_2_tdata2[30] == dec_i0_match_data_2[30]; // @[el2_lib.scala 219:79]
  wire  _T_893 = _T_889 | _T_892; // @[el2_lib.scala 219:24]
  wire  _T_895 = &io_trigger_pkt_any_2_tdata2[30:0]; // @[el2_lib.scala 219:37]
  wire  _T_896 = _T_895 & _T_679; // @[el2_lib.scala 219:42]
  wire  _T_899 = io_trigger_pkt_any_2_tdata2[31] == dec_i0_match_data_2[31]; // @[el2_lib.scala 219:79]
  wire  _T_900 = _T_896 | _T_899; // @[el2_lib.scala 219:24]
  wire [7:0] _T_907 = {_T_732,_T_725,_T_718,_T_711,_T_704,_T_697,_T_690,_T_683}; // @[el2_lib.scala 220:14]
  wire [15:0] _T_915 = {_T_788,_T_781,_T_774,_T_767,_T_760,_T_753,_T_746,_T_739,_T_907}; // @[el2_lib.scala 220:14]
  wire [7:0] _T_922 = {_T_844,_T_837,_T_830,_T_823,_T_816,_T_809,_T_802,_T_795}; // @[el2_lib.scala 220:14]
  wire [31:0] _T_931 = {_T_900,_T_893,_T_886,_T_879,_T_872,_T_865,_T_858,_T_851,_T_922,_T_915}; // @[el2_lib.scala 220:14]
  wire  _T_932 = &_T_931; // @[el2_lib.scala 220:21]
  wire  _T_933 = _T_672 & _T_932; // @[el2_dec_trigger.scala 15:109]
  wire  _T_934 = io_trigger_pkt_any_3_execute & io_trigger_pkt_any_3_m; // @[el2_dec_trigger.scala 15:83]
  wire  _T_939 = &io_trigger_pkt_any_3_tdata2; // @[el2_lib.scala 216:73]
  wire  _T_940 = ~_T_939; // @[el2_lib.scala 216:47]
  wire  _T_941 = io_trigger_pkt_any_3_match_ & _T_940; // @[el2_lib.scala 216:44]
  wire  _T_944 = io_trigger_pkt_any_3_tdata2[0] == dec_i0_match_data_3[0]; // @[el2_lib.scala 217:52]
  wire  _T_945 = _T_941 | _T_944; // @[el2_lib.scala 217:41]
  wire  _T_947 = &io_trigger_pkt_any_3_tdata2[0]; // @[el2_lib.scala 219:37]
  wire  _T_948 = _T_947 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_951 = io_trigger_pkt_any_3_tdata2[1] == dec_i0_match_data_3[1]; // @[el2_lib.scala 219:79]
  wire  _T_952 = _T_948 | _T_951; // @[el2_lib.scala 219:24]
  wire  _T_954 = &io_trigger_pkt_any_3_tdata2[1:0]; // @[el2_lib.scala 219:37]
  wire  _T_955 = _T_954 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_958 = io_trigger_pkt_any_3_tdata2[2] == dec_i0_match_data_3[2]; // @[el2_lib.scala 219:79]
  wire  _T_959 = _T_955 | _T_958; // @[el2_lib.scala 219:24]
  wire  _T_961 = &io_trigger_pkt_any_3_tdata2[2:0]; // @[el2_lib.scala 219:37]
  wire  _T_962 = _T_961 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_965 = io_trigger_pkt_any_3_tdata2[3] == dec_i0_match_data_3[3]; // @[el2_lib.scala 219:79]
  wire  _T_966 = _T_962 | _T_965; // @[el2_lib.scala 219:24]
  wire  _T_968 = &io_trigger_pkt_any_3_tdata2[3:0]; // @[el2_lib.scala 219:37]
  wire  _T_969 = _T_968 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_972 = io_trigger_pkt_any_3_tdata2[4] == dec_i0_match_data_3[4]; // @[el2_lib.scala 219:79]
  wire  _T_973 = _T_969 | _T_972; // @[el2_lib.scala 219:24]
  wire  _T_975 = &io_trigger_pkt_any_3_tdata2[4:0]; // @[el2_lib.scala 219:37]
  wire  _T_976 = _T_975 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_979 = io_trigger_pkt_any_3_tdata2[5] == dec_i0_match_data_3[5]; // @[el2_lib.scala 219:79]
  wire  _T_980 = _T_976 | _T_979; // @[el2_lib.scala 219:24]
  wire  _T_982 = &io_trigger_pkt_any_3_tdata2[5:0]; // @[el2_lib.scala 219:37]
  wire  _T_983 = _T_982 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_986 = io_trigger_pkt_any_3_tdata2[6] == dec_i0_match_data_3[6]; // @[el2_lib.scala 219:79]
  wire  _T_987 = _T_983 | _T_986; // @[el2_lib.scala 219:24]
  wire  _T_989 = &io_trigger_pkt_any_3_tdata2[6:0]; // @[el2_lib.scala 219:37]
  wire  _T_990 = _T_989 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_993 = io_trigger_pkt_any_3_tdata2[7] == dec_i0_match_data_3[7]; // @[el2_lib.scala 219:79]
  wire  _T_994 = _T_990 | _T_993; // @[el2_lib.scala 219:24]
  wire  _T_996 = &io_trigger_pkt_any_3_tdata2[7:0]; // @[el2_lib.scala 219:37]
  wire  _T_997 = _T_996 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1000 = io_trigger_pkt_any_3_tdata2[8] == dec_i0_match_data_3[8]; // @[el2_lib.scala 219:79]
  wire  _T_1001 = _T_997 | _T_1000; // @[el2_lib.scala 219:24]
  wire  _T_1003 = &io_trigger_pkt_any_3_tdata2[8:0]; // @[el2_lib.scala 219:37]
  wire  _T_1004 = _T_1003 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1007 = io_trigger_pkt_any_3_tdata2[9] == dec_i0_match_data_3[9]; // @[el2_lib.scala 219:79]
  wire  _T_1008 = _T_1004 | _T_1007; // @[el2_lib.scala 219:24]
  wire  _T_1010 = &io_trigger_pkt_any_3_tdata2[9:0]; // @[el2_lib.scala 219:37]
  wire  _T_1011 = _T_1010 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1014 = io_trigger_pkt_any_3_tdata2[10] == dec_i0_match_data_3[10]; // @[el2_lib.scala 219:79]
  wire  _T_1015 = _T_1011 | _T_1014; // @[el2_lib.scala 219:24]
  wire  _T_1017 = &io_trigger_pkt_any_3_tdata2[10:0]; // @[el2_lib.scala 219:37]
  wire  _T_1018 = _T_1017 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1021 = io_trigger_pkt_any_3_tdata2[11] == dec_i0_match_data_3[11]; // @[el2_lib.scala 219:79]
  wire  _T_1022 = _T_1018 | _T_1021; // @[el2_lib.scala 219:24]
  wire  _T_1024 = &io_trigger_pkt_any_3_tdata2[11:0]; // @[el2_lib.scala 219:37]
  wire  _T_1025 = _T_1024 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1028 = io_trigger_pkt_any_3_tdata2[12] == dec_i0_match_data_3[12]; // @[el2_lib.scala 219:79]
  wire  _T_1029 = _T_1025 | _T_1028; // @[el2_lib.scala 219:24]
  wire  _T_1031 = &io_trigger_pkt_any_3_tdata2[12:0]; // @[el2_lib.scala 219:37]
  wire  _T_1032 = _T_1031 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1035 = io_trigger_pkt_any_3_tdata2[13] == dec_i0_match_data_3[13]; // @[el2_lib.scala 219:79]
  wire  _T_1036 = _T_1032 | _T_1035; // @[el2_lib.scala 219:24]
  wire  _T_1038 = &io_trigger_pkt_any_3_tdata2[13:0]; // @[el2_lib.scala 219:37]
  wire  _T_1039 = _T_1038 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1042 = io_trigger_pkt_any_3_tdata2[14] == dec_i0_match_data_3[14]; // @[el2_lib.scala 219:79]
  wire  _T_1043 = _T_1039 | _T_1042; // @[el2_lib.scala 219:24]
  wire  _T_1045 = &io_trigger_pkt_any_3_tdata2[14:0]; // @[el2_lib.scala 219:37]
  wire  _T_1046 = _T_1045 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1049 = io_trigger_pkt_any_3_tdata2[15] == dec_i0_match_data_3[15]; // @[el2_lib.scala 219:79]
  wire  _T_1050 = _T_1046 | _T_1049; // @[el2_lib.scala 219:24]
  wire  _T_1052 = &io_trigger_pkt_any_3_tdata2[15:0]; // @[el2_lib.scala 219:37]
  wire  _T_1053 = _T_1052 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1056 = io_trigger_pkt_any_3_tdata2[16] == dec_i0_match_data_3[16]; // @[el2_lib.scala 219:79]
  wire  _T_1057 = _T_1053 | _T_1056; // @[el2_lib.scala 219:24]
  wire  _T_1059 = &io_trigger_pkt_any_3_tdata2[16:0]; // @[el2_lib.scala 219:37]
  wire  _T_1060 = _T_1059 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1063 = io_trigger_pkt_any_3_tdata2[17] == dec_i0_match_data_3[17]; // @[el2_lib.scala 219:79]
  wire  _T_1064 = _T_1060 | _T_1063; // @[el2_lib.scala 219:24]
  wire  _T_1066 = &io_trigger_pkt_any_3_tdata2[17:0]; // @[el2_lib.scala 219:37]
  wire  _T_1067 = _T_1066 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1070 = io_trigger_pkt_any_3_tdata2[18] == dec_i0_match_data_3[18]; // @[el2_lib.scala 219:79]
  wire  _T_1071 = _T_1067 | _T_1070; // @[el2_lib.scala 219:24]
  wire  _T_1073 = &io_trigger_pkt_any_3_tdata2[18:0]; // @[el2_lib.scala 219:37]
  wire  _T_1074 = _T_1073 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1077 = io_trigger_pkt_any_3_tdata2[19] == dec_i0_match_data_3[19]; // @[el2_lib.scala 219:79]
  wire  _T_1078 = _T_1074 | _T_1077; // @[el2_lib.scala 219:24]
  wire  _T_1080 = &io_trigger_pkt_any_3_tdata2[19:0]; // @[el2_lib.scala 219:37]
  wire  _T_1081 = _T_1080 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1084 = io_trigger_pkt_any_3_tdata2[20] == dec_i0_match_data_3[20]; // @[el2_lib.scala 219:79]
  wire  _T_1085 = _T_1081 | _T_1084; // @[el2_lib.scala 219:24]
  wire  _T_1087 = &io_trigger_pkt_any_3_tdata2[20:0]; // @[el2_lib.scala 219:37]
  wire  _T_1088 = _T_1087 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1091 = io_trigger_pkt_any_3_tdata2[21] == dec_i0_match_data_3[21]; // @[el2_lib.scala 219:79]
  wire  _T_1092 = _T_1088 | _T_1091; // @[el2_lib.scala 219:24]
  wire  _T_1094 = &io_trigger_pkt_any_3_tdata2[21:0]; // @[el2_lib.scala 219:37]
  wire  _T_1095 = _T_1094 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1098 = io_trigger_pkt_any_3_tdata2[22] == dec_i0_match_data_3[22]; // @[el2_lib.scala 219:79]
  wire  _T_1099 = _T_1095 | _T_1098; // @[el2_lib.scala 219:24]
  wire  _T_1101 = &io_trigger_pkt_any_3_tdata2[22:0]; // @[el2_lib.scala 219:37]
  wire  _T_1102 = _T_1101 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1105 = io_trigger_pkt_any_3_tdata2[23] == dec_i0_match_data_3[23]; // @[el2_lib.scala 219:79]
  wire  _T_1106 = _T_1102 | _T_1105; // @[el2_lib.scala 219:24]
  wire  _T_1108 = &io_trigger_pkt_any_3_tdata2[23:0]; // @[el2_lib.scala 219:37]
  wire  _T_1109 = _T_1108 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1112 = io_trigger_pkt_any_3_tdata2[24] == dec_i0_match_data_3[24]; // @[el2_lib.scala 219:79]
  wire  _T_1113 = _T_1109 | _T_1112; // @[el2_lib.scala 219:24]
  wire  _T_1115 = &io_trigger_pkt_any_3_tdata2[24:0]; // @[el2_lib.scala 219:37]
  wire  _T_1116 = _T_1115 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1119 = io_trigger_pkt_any_3_tdata2[25] == dec_i0_match_data_3[25]; // @[el2_lib.scala 219:79]
  wire  _T_1120 = _T_1116 | _T_1119; // @[el2_lib.scala 219:24]
  wire  _T_1122 = &io_trigger_pkt_any_3_tdata2[25:0]; // @[el2_lib.scala 219:37]
  wire  _T_1123 = _T_1122 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1126 = io_trigger_pkt_any_3_tdata2[26] == dec_i0_match_data_3[26]; // @[el2_lib.scala 219:79]
  wire  _T_1127 = _T_1123 | _T_1126; // @[el2_lib.scala 219:24]
  wire  _T_1129 = &io_trigger_pkt_any_3_tdata2[26:0]; // @[el2_lib.scala 219:37]
  wire  _T_1130 = _T_1129 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1133 = io_trigger_pkt_any_3_tdata2[27] == dec_i0_match_data_3[27]; // @[el2_lib.scala 219:79]
  wire  _T_1134 = _T_1130 | _T_1133; // @[el2_lib.scala 219:24]
  wire  _T_1136 = &io_trigger_pkt_any_3_tdata2[27:0]; // @[el2_lib.scala 219:37]
  wire  _T_1137 = _T_1136 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1140 = io_trigger_pkt_any_3_tdata2[28] == dec_i0_match_data_3[28]; // @[el2_lib.scala 219:79]
  wire  _T_1141 = _T_1137 | _T_1140; // @[el2_lib.scala 219:24]
  wire  _T_1143 = &io_trigger_pkt_any_3_tdata2[28:0]; // @[el2_lib.scala 219:37]
  wire  _T_1144 = _T_1143 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1147 = io_trigger_pkt_any_3_tdata2[29] == dec_i0_match_data_3[29]; // @[el2_lib.scala 219:79]
  wire  _T_1148 = _T_1144 | _T_1147; // @[el2_lib.scala 219:24]
  wire  _T_1150 = &io_trigger_pkt_any_3_tdata2[29:0]; // @[el2_lib.scala 219:37]
  wire  _T_1151 = _T_1150 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1154 = io_trigger_pkt_any_3_tdata2[30] == dec_i0_match_data_3[30]; // @[el2_lib.scala 219:79]
  wire  _T_1155 = _T_1151 | _T_1154; // @[el2_lib.scala 219:24]
  wire  _T_1157 = &io_trigger_pkt_any_3_tdata2[30:0]; // @[el2_lib.scala 219:37]
  wire  _T_1158 = _T_1157 & _T_941; // @[el2_lib.scala 219:42]
  wire  _T_1161 = io_trigger_pkt_any_3_tdata2[31] == dec_i0_match_data_3[31]; // @[el2_lib.scala 219:79]
  wire  _T_1162 = _T_1158 | _T_1161; // @[el2_lib.scala 219:24]
  wire [7:0] _T_1169 = {_T_994,_T_987,_T_980,_T_973,_T_966,_T_959,_T_952,_T_945}; // @[el2_lib.scala 220:14]
  wire [15:0] _T_1177 = {_T_1050,_T_1043,_T_1036,_T_1029,_T_1022,_T_1015,_T_1008,_T_1001,_T_1169}; // @[el2_lib.scala 220:14]
  wire [7:0] _T_1184 = {_T_1106,_T_1099,_T_1092,_T_1085,_T_1078,_T_1071,_T_1064,_T_1057}; // @[el2_lib.scala 220:14]
  wire [31:0] _T_1193 = {_T_1162,_T_1155,_T_1148,_T_1141,_T_1134,_T_1127,_T_1120,_T_1113,_T_1184,_T_1177}; // @[el2_lib.scala 220:14]
  wire  _T_1194 = &_T_1193; // @[el2_lib.scala 220:21]
  wire  _T_1195 = _T_934 & _T_1194; // @[el2_dec_trigger.scala 15:109]
  wire [2:0] _T_1197 = {_T_1195,_T_933,_T_671}; // @[Cat.scala 29:58]
  assign io_dec_i0_trigger_match_d = {_T_1197,_T_409}; // @[el2_dec_trigger.scala 15:29]
endmodule
