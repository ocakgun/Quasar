module rvclkhdr(
  output  io_l1clk,
  input   io_clk,
  input   io_en,
  input   io_scan_mode
);
  wire  clkhdr_Q; // @[el2_lib.scala 474:26]
  wire  clkhdr_CK; // @[el2_lib.scala 474:26]
  wire  clkhdr_EN; // @[el2_lib.scala 474:26]
  wire  clkhdr_SE; // @[el2_lib.scala 474:26]
  gated_latch clkhdr ( // @[el2_lib.scala 474:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign io_l1clk = clkhdr_Q; // @[el2_lib.scala 475:14]
  assign clkhdr_CK = io_clk; // @[el2_lib.scala 476:18]
  assign clkhdr_EN = io_en; // @[el2_lib.scala 477:18]
  assign clkhdr_SE = io_scan_mode; // @[el2_lib.scala 478:18]
endmodule
module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [95:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [63:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [63:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_1_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_2_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_3_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_4_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_5_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_6_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_7_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_8_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_9_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_10_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_11_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_12_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_13_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_14_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_15_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_16_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_17_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_18_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_19_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_20_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_21_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_22_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_23_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_24_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_25_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_26_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_27_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_28_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_29_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_30_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_31_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_32_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_33_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_34_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_35_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_36_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_37_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_38_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_39_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_40_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_41_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_42_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_43_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_44_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_45_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_46_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_47_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_48_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_49_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_50_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_51_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_52_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_53_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_54_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_55_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_56_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_57_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_58_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_59_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_60_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_61_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_62_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_63_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_64_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_65_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_66_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_67_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_68_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_69_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_70_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_71_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_72_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_73_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_74_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_75_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_76_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_77_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_78_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_79_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_80_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_81_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_82_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_83_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_84_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_85_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_86_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_87_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_88_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_89_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_90_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_91_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_92_io_scan_mode; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_l1clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_clk; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_en; // @[el2_lib.scala 483:22]
  wire  rvclkhdr_93_io_scan_mode; // @[el2_lib.scala 483:22]
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 186:53]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 322:61]
  wire  _T_319 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 323:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_319; // @[el2_ifu_mem_ctl.scala 323:42]
  wire  _T = io_ifc_fetch_req_bf_raw | ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 187:53]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 254:30]
  wire  _T_1 = _T | miss_pending; // @[el2_ifu_mem_ctl.scala 187:71]
  wire  _T_2 = _T_1 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 187:86]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 557:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_319; // @[el2_ifu_mem_ctl.scala 559:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 188:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 309:63]
  wire [4:0] _GEN_436 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 675:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_436 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 675:53]
  wire  _T_3128 = |ic_fetch_val_shift_right[3:2]; // @[el2_ifu_mem_ctl.scala 678:91]
  wire  _T_3130 = _T_3128 & _T_319; // @[el2_ifu_mem_ctl.scala 678:95]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 324:60]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 276:46]
  wire  _T_3131 = _T_3130 & fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 678:117]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 664:59]
  wire  _T_3132 = _T_3131 | iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 678:134]
  wire  _T_3133 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 678:158]
  wire  _T_3134 = _T_3132 & _T_3133; // @[el2_ifu_mem_ctl.scala 678:156]
  wire  _T_3120 = |ic_fetch_val_shift_right[1:0]; // @[el2_ifu_mem_ctl.scala 678:91]
  wire  _T_3122 = _T_3120 & _T_319; // @[el2_ifu_mem_ctl.scala 678:95]
  wire  _T_3123 = _T_3122 & fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 678:117]
  wire  _T_3124 = _T_3123 | iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 678:134]
  wire  _T_3126 = _T_3124 & _T_3133; // @[el2_ifu_mem_ctl.scala 678:156]
  wire [1:0] iccm_ecc_word_enable = {_T_3134,_T_3126}; // @[Cat.scala 29:58]
  wire  _T_3234 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 333:30]
  wire  _T_3235 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 333:44]
  wire  _T_3236 = _T_3234 ^ _T_3235; // @[el2_lib.scala 333:35]
  wire [5:0] _T_3244 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 333:76]
  wire  _T_3245 = ^_T_3244; // @[el2_lib.scala 333:83]
  wire  _T_3246 = io_iccm_rd_data_ecc[37] ^ _T_3245; // @[el2_lib.scala 333:71]
  wire [6:0] _T_3253 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 333:103]
  wire [14:0] _T_3261 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3253}; // @[el2_lib.scala 333:103]
  wire  _T_3262 = ^_T_3261; // @[el2_lib.scala 333:110]
  wire  _T_3263 = io_iccm_rd_data_ecc[36] ^ _T_3262; // @[el2_lib.scala 333:98]
  wire [6:0] _T_3270 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 333:130]
  wire [14:0] _T_3278 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3270}; // @[el2_lib.scala 333:130]
  wire  _T_3279 = ^_T_3278; // @[el2_lib.scala 333:137]
  wire  _T_3280 = io_iccm_rd_data_ecc[35] ^ _T_3279; // @[el2_lib.scala 333:125]
  wire [8:0] _T_3289 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 333:157]
  wire [17:0] _T_3298 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3289}; // @[el2_lib.scala 333:157]
  wire  _T_3299 = ^_T_3298; // @[el2_lib.scala 333:164]
  wire  _T_3300 = io_iccm_rd_data_ecc[34] ^ _T_3299; // @[el2_lib.scala 333:152]
  wire [8:0] _T_3309 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 333:184]
  wire [17:0] _T_3318 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3309}; // @[el2_lib.scala 333:184]
  wire  _T_3319 = ^_T_3318; // @[el2_lib.scala 333:191]
  wire  _T_3320 = io_iccm_rd_data_ecc[33] ^ _T_3319; // @[el2_lib.scala 333:179]
  wire [8:0] _T_3329 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 333:211]
  wire [17:0] _T_3338 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3329}; // @[el2_lib.scala 333:211]
  wire  _T_3339 = ^_T_3338; // @[el2_lib.scala 333:218]
  wire  _T_3340 = io_iccm_rd_data_ecc[32] ^ _T_3339; // @[el2_lib.scala 333:206]
  wire [6:0] _T_3346 = {_T_3236,_T_3246,_T_3263,_T_3280,_T_3300,_T_3320,_T_3340}; // @[Cat.scala 29:58]
  wire  _T_3347 = _T_3346 != 7'h0; // @[el2_lib.scala 334:44]
  wire  _T_3348 = iccm_ecc_word_enable[0] & _T_3347; // @[el2_lib.scala 334:32]
  wire  _T_3350 = _T_3348 & _T_3346[6]; // @[el2_lib.scala 334:53]
  wire  _T_3619 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 333:30]
  wire  _T_3620 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 333:44]
  wire  _T_3621 = _T_3619 ^ _T_3620; // @[el2_lib.scala 333:35]
  wire [5:0] _T_3629 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 333:76]
  wire  _T_3630 = ^_T_3629; // @[el2_lib.scala 333:83]
  wire  _T_3631 = io_iccm_rd_data_ecc[76] ^ _T_3630; // @[el2_lib.scala 333:71]
  wire [6:0] _T_3638 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 333:103]
  wire [14:0] _T_3646 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3638}; // @[el2_lib.scala 333:103]
  wire  _T_3647 = ^_T_3646; // @[el2_lib.scala 333:110]
  wire  _T_3648 = io_iccm_rd_data_ecc[75] ^ _T_3647; // @[el2_lib.scala 333:98]
  wire [6:0] _T_3655 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 333:130]
  wire [14:0] _T_3663 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3655}; // @[el2_lib.scala 333:130]
  wire  _T_3664 = ^_T_3663; // @[el2_lib.scala 333:137]
  wire  _T_3665 = io_iccm_rd_data_ecc[74] ^ _T_3664; // @[el2_lib.scala 333:125]
  wire [8:0] _T_3674 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 333:157]
  wire [17:0] _T_3683 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3674}; // @[el2_lib.scala 333:157]
  wire  _T_3684 = ^_T_3683; // @[el2_lib.scala 333:164]
  wire  _T_3685 = io_iccm_rd_data_ecc[73] ^ _T_3684; // @[el2_lib.scala 333:152]
  wire [8:0] _T_3694 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 333:184]
  wire [17:0] _T_3703 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3694}; // @[el2_lib.scala 333:184]
  wire  _T_3704 = ^_T_3703; // @[el2_lib.scala 333:191]
  wire  _T_3705 = io_iccm_rd_data_ecc[72] ^ _T_3704; // @[el2_lib.scala 333:179]
  wire [8:0] _T_3714 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 333:211]
  wire [17:0] _T_3723 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3714}; // @[el2_lib.scala 333:211]
  wire  _T_3724 = ^_T_3723; // @[el2_lib.scala 333:218]
  wire  _T_3725 = io_iccm_rd_data_ecc[71] ^ _T_3724; // @[el2_lib.scala 333:206]
  wire [6:0] _T_3731 = {_T_3621,_T_3631,_T_3648,_T_3665,_T_3685,_T_3705,_T_3725}; // @[Cat.scala 29:58]
  wire  _T_3732 = _T_3731 != 7'h0; // @[el2_lib.scala 334:44]
  wire  _T_3733 = iccm_ecc_word_enable[1] & _T_3732; // @[el2_lib.scala 334:32]
  wire  _T_3735 = _T_3733 & _T_3731[6]; // @[el2_lib.scala 334:53]
  wire [1:0] iccm_single_ecc_error = {_T_3350,_T_3735}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 191:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 641:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 192:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 193:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 484:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 193:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 193:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 193:72]
  wire  _T_2525 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2530 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2550 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 534:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 398:42]
  wire  _T_2552 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 534:79]
  wire  _T_2553 = _T_2550 | _T_2552; // @[el2_ifu_mem_ctl.scala 534:56]
  wire  _T_2554 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 534:122]
  wire  _T_2555 = ~_T_2554; // @[el2_ifu_mem_ctl.scala 534:101]
  wire  _T_2556 = _T_2553 & _T_2555; // @[el2_ifu_mem_ctl.scala 534:99]
  wire  _T_2557 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2571 = io_ifu_fetch_val[0] & _T_319; // @[el2_ifu_mem_ctl.scala 541:45]
  wire  _T_2572 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 541:69]
  wire  _T_2573 = _T_2571 & _T_2572; // @[el2_ifu_mem_ctl.scala 541:67]
  wire  _T_2574 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_37 = _T_2557 ? _T_2573 : _T_2574; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_2530 ? _T_2556 : _GEN_37; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2525 ? 1'h0 : _GEN_41; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 193:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 195:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 195:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 284:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 284:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 710:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 284:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 275:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 275:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 326:71]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 275:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 275:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 284:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 284:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 284:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 284:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 284:114]
  reg  ifu_bus_rvalid_unq_ff; // @[el2_ifu_mem_ctl.scala 584:56]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 556:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 598:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 625:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 311:62]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 606:56]
  wire  _T_2671 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 623:69]
  wire  _T_2672 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 623:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2671 : _T_2672; // @[el2_ifu_mem_ctl.scala 623:28]
  wire  _T_2623 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 602:68]
  wire  _T_2624 = ic_act_miss_f | _T_2623; // @[el2_ifu_mem_ctl.scala 602:48]
  wire  bus_reset_data_beat_cnt = _T_2624 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 602:91]
  wire  _T_2620 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 601:50]
  wire  _T_2621 = bus_ifu_wr_en_ff & _T_2620; // @[el2_ifu_mem_ctl.scala 601:48]
  wire  _T_2622 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 601:72]
  wire  bus_inc_data_beat_cnt = _T_2621 & _T_2622; // @[el2_ifu_mem_ctl.scala 601:70]
  wire [2:0] _T_2628 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 605:115]
  wire [2:0] _T_2630 = bus_inc_data_beat_cnt ? _T_2628 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2625 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 603:32]
  wire  _T_2626 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 603:57]
  wire  bus_hold_data_beat_cnt = _T_2625 & _T_2626; // @[el2_ifu_mem_ctl.scala 603:55]
  wire [2:0] _T_2631 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2630 | _T_2631; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 195:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 195:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 196:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 195:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 196:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_319; // @[el2_ifu_mem_ctl.scala 202:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 202:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 435:45]
  wire  _T_2154 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 457:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 412:60]
  wire  _T_2185 = _T_2154 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2158 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 457:127]
  wire  _T_2186 = _T_2158 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2193 = _T_2185 | _T_2186; // @[Mux.scala 27:72]
  wire  _T_2162 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 457:127]
  wire  _T_2187 = _T_2162 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2194 = _T_2193 | _T_2187; // @[Mux.scala 27:72]
  wire  _T_2166 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 457:127]
  wire  _T_2188 = _T_2166 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2195 = _T_2194 | _T_2188; // @[Mux.scala 27:72]
  wire  _T_2170 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 457:127]
  wire  _T_2189 = _T_2170 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2196 = _T_2195 | _T_2189; // @[Mux.scala 27:72]
  wire  _T_2174 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 457:127]
  wire  _T_2190 = _T_2174 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2197 = _T_2196 | _T_2190; // @[Mux.scala 27:72]
  wire  _T_2178 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 457:127]
  wire  _T_2191 = _T_2178 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2198 = _T_2197 | _T_2191; // @[Mux.scala 27:72]
  wire  _T_2182 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 457:127]
  wire  _T_2192 = _T_2182 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2198 | _T_2192; // @[Mux.scala 27:72]
  wire  _T_2240 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 459:69]
  wire  _T_2241 = ic_miss_buff_data_valid_bypass_index & _T_2240; // @[el2_ifu_mem_ctl.scala 459:67]
  wire  _T_2243 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 459:91]
  wire  _T_2244 = _T_2241 & _T_2243; // @[el2_ifu_mem_ctl.scala 459:89]
  wire  _T_2249 = _T_2241 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 460:65]
  wire  _T_2250 = _T_2244 | _T_2249; // @[el2_ifu_mem_ctl.scala 459:112]
  wire  _T_2252 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 461:43]
  wire  _T_2255 = _T_2252 & _T_2243; // @[el2_ifu_mem_ctl.scala 461:65]
  wire  _T_2256 = _T_2250 | _T_2255; // @[el2_ifu_mem_ctl.scala 460:88]
  wire  _T_2260 = _T_2252 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 462:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 438:75]
  wire  _T_2200 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 458:110]
  wire  _T_2224 = _T_2200 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2203 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 458:110]
  wire  _T_2225 = _T_2203 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2232 = _T_2224 | _T_2225; // @[Mux.scala 27:72]
  wire  _T_2206 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 458:110]
  wire  _T_2226 = _T_2206 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2233 = _T_2232 | _T_2226; // @[Mux.scala 27:72]
  wire  _T_2209 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 458:110]
  wire  _T_2227 = _T_2209 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2234 = _T_2233 | _T_2227; // @[Mux.scala 27:72]
  wire  _T_2212 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 458:110]
  wire  _T_2228 = _T_2212 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2235 = _T_2234 | _T_2228; // @[Mux.scala 27:72]
  wire  _T_2215 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 458:110]
  wire  _T_2229 = _T_2215 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2236 = _T_2235 | _T_2229; // @[Mux.scala 27:72]
  wire  _T_2218 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 458:110]
  wire  _T_2230 = _T_2218 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2237 = _T_2236 | _T_2230; // @[Mux.scala 27:72]
  wire  _T_2221 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 458:110]
  wire  _T_2231 = _T_2221 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2237 | _T_2231; // @[Mux.scala 27:72]
  wire  _T_2261 = _T_2260 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 462:87]
  wire  _T_2262 = _T_2256 | _T_2261; // @[el2_ifu_mem_ctl.scala 461:88]
  wire  _T_2266 = ic_miss_buff_data_valid_bypass_index & _T_2182; // @[el2_ifu_mem_ctl.scala 463:43]
  wire  miss_buff_hit_unq_f = _T_2262 | _T_2266; // @[el2_ifu_mem_ctl.scala 462:131]
  wire  _T_2282 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 468:55]
  wire  _T_2283 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 468:87]
  wire  _T_2284 = _T_2282 | _T_2283; // @[el2_ifu_mem_ctl.scala 468:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2284; // @[el2_ifu_mem_ctl.scala 468:41]
  wire  _T_2267 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 465:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 312:49]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[el2_ifu_mem_ctl.scala 456:51]
  wire  _T_2268 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 465:68]
  wire  _T_2269 = miss_buff_hit_unq_f & _T_2268; // @[el2_ifu_mem_ctl.scala 465:66]
  wire  stream_hit_f = _T_2267 & _T_2269; // @[el2_ifu_mem_ctl.scala 465:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 279:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 279:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 279:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 608:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 635:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 206:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 206:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 206:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 206:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 206:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 207:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 207:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 207:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 208:16]
  wire  _T_44 = _T_42 & _T_319; // @[el2_ifu_mem_ctl.scala 208:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 208:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 208:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 209:49]
  wire  _T_54 = ic_byp_hit_f & _T_319; // @[el2_ifu_mem_ctl.scala 210:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 210:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 210:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 198:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 210:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 210:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 210:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_319; // @[el2_ifu_mem_ctl.scala 211:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 211:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 211:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 211:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 212:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 213:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 213:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 213:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 212:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 211:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 210:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 209:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 208:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 207:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 206:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2279 = byp_fetch_index[4:1] == 4'hf; // @[el2_ifu_mem_ctl.scala 467:60]
  wire  _T_2280 = _T_2279 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 467:94]
  wire  stream_eol_f = _T_2280 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 467:112]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 221:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 221:87]
  wire  _T_113 = _T_111 & _T_2622; // @[el2_ifu_mem_ctl.scala 221:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 221:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 225:48]
  wire  _T_126 = _T_124 & _T_2622; // @[el2_ifu_mem_ctl.scala 225:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 225:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 285:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 285:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 285:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 285:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 285:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 286:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 285:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 286:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 340:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 286:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 286:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 286:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 229:50]
  wire  _T_137 = _T_135 & _T_2622; // @[el2_ifu_mem_ctl.scala 229:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 287:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 288:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 288:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 287:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 230:35]
  wire  _T_143 = _T_141 & _T_2622; // @[el2_ifu_mem_ctl.scala 230:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 230:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 229:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 235:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 234:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 234:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 239:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 239:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 196:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 196:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 196:26]
  wire  _T_30 = ic_act_miss_f & _T_2622; // @[el2_ifu_mem_ctl.scala 203:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 214:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 214:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 214:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 214:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 214:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 214:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 218:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 218:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 218:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 222:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 222:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 226:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 226:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 231:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 231:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 231:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 236:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 236:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 255:95]
  wire  _T_175 = _T_2282 & _T_174; // @[el2_ifu_mem_ctl.scala 255:93]
  wire  crit_wd_byp_ok_ff = _T_2283 | _T_175; // @[el2_ifu_mem_ctl.scala 255:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 256:36]
  wire  _T_180 = _T_2282 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 256:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 256:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 256:70]
  wire  _T_184 = _T_2282 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 257:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 257:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 256:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 257:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 258:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 258:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 257:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 260:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 260:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:64]
  reg [6:0] ifu_ic_rw_int_addr_ff; // @[el2_ifu_mem_ctl.scala 742:14]
  wire  _T_4670 = ifu_ic_rw_int_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_0; // @[Reg.scala 27:20]
  wire  _T_4798 = _T_4670 & way_status_out_0; // @[Mux.scala 27:72]
  wire  _T_4671 = ifu_ic_rw_int_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_1; // @[Reg.scala 27:20]
  wire  _T_4799 = _T_4671 & way_status_out_1; // @[Mux.scala 27:72]
  wire  _T_4926 = _T_4798 | _T_4799; // @[Mux.scala 27:72]
  wire  _T_4672 = ifu_ic_rw_int_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_2; // @[Reg.scala 27:20]
  wire  _T_4800 = _T_4672 & way_status_out_2; // @[Mux.scala 27:72]
  wire  _T_4927 = _T_4926 | _T_4800; // @[Mux.scala 27:72]
  wire  _T_4673 = ifu_ic_rw_int_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_3; // @[Reg.scala 27:20]
  wire  _T_4801 = _T_4673 & way_status_out_3; // @[Mux.scala 27:72]
  wire  _T_4928 = _T_4927 | _T_4801; // @[Mux.scala 27:72]
  wire  _T_4674 = ifu_ic_rw_int_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_4; // @[Reg.scala 27:20]
  wire  _T_4802 = _T_4674 & way_status_out_4; // @[Mux.scala 27:72]
  wire  _T_4929 = _T_4928 | _T_4802; // @[Mux.scala 27:72]
  wire  _T_4675 = ifu_ic_rw_int_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_5; // @[Reg.scala 27:20]
  wire  _T_4803 = _T_4675 & way_status_out_5; // @[Mux.scala 27:72]
  wire  _T_4930 = _T_4929 | _T_4803; // @[Mux.scala 27:72]
  wire  _T_4676 = ifu_ic_rw_int_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_6; // @[Reg.scala 27:20]
  wire  _T_4804 = _T_4676 & way_status_out_6; // @[Mux.scala 27:72]
  wire  _T_4931 = _T_4930 | _T_4804; // @[Mux.scala 27:72]
  wire  _T_4677 = ifu_ic_rw_int_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_7; // @[Reg.scala 27:20]
  wire  _T_4805 = _T_4677 & way_status_out_7; // @[Mux.scala 27:72]
  wire  _T_4932 = _T_4931 | _T_4805; // @[Mux.scala 27:72]
  wire  _T_4678 = ifu_ic_rw_int_addr_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_8; // @[Reg.scala 27:20]
  wire  _T_4806 = _T_4678 & way_status_out_8; // @[Mux.scala 27:72]
  wire  _T_4933 = _T_4932 | _T_4806; // @[Mux.scala 27:72]
  wire  _T_4679 = ifu_ic_rw_int_addr_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_9; // @[Reg.scala 27:20]
  wire  _T_4807 = _T_4679 & way_status_out_9; // @[Mux.scala 27:72]
  wire  _T_4934 = _T_4933 | _T_4807; // @[Mux.scala 27:72]
  wire  _T_4680 = ifu_ic_rw_int_addr_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_10; // @[Reg.scala 27:20]
  wire  _T_4808 = _T_4680 & way_status_out_10; // @[Mux.scala 27:72]
  wire  _T_4935 = _T_4934 | _T_4808; // @[Mux.scala 27:72]
  wire  _T_4681 = ifu_ic_rw_int_addr_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_11; // @[Reg.scala 27:20]
  wire  _T_4809 = _T_4681 & way_status_out_11; // @[Mux.scala 27:72]
  wire  _T_4936 = _T_4935 | _T_4809; // @[Mux.scala 27:72]
  wire  _T_4682 = ifu_ic_rw_int_addr_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_12; // @[Reg.scala 27:20]
  wire  _T_4810 = _T_4682 & way_status_out_12; // @[Mux.scala 27:72]
  wire  _T_4937 = _T_4936 | _T_4810; // @[Mux.scala 27:72]
  wire  _T_4683 = ifu_ic_rw_int_addr_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_13; // @[Reg.scala 27:20]
  wire  _T_4811 = _T_4683 & way_status_out_13; // @[Mux.scala 27:72]
  wire  _T_4938 = _T_4937 | _T_4811; // @[Mux.scala 27:72]
  wire  _T_4684 = ifu_ic_rw_int_addr_ff == 7'he; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_14; // @[Reg.scala 27:20]
  wire  _T_4812 = _T_4684 & way_status_out_14; // @[Mux.scala 27:72]
  wire  _T_4939 = _T_4938 | _T_4812; // @[Mux.scala 27:72]
  wire  _T_4685 = ifu_ic_rw_int_addr_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_15; // @[Reg.scala 27:20]
  wire  _T_4813 = _T_4685 & way_status_out_15; // @[Mux.scala 27:72]
  wire  _T_4940 = _T_4939 | _T_4813; // @[Mux.scala 27:72]
  wire  _T_4686 = ifu_ic_rw_int_addr_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_16; // @[Reg.scala 27:20]
  wire  _T_4814 = _T_4686 & way_status_out_16; // @[Mux.scala 27:72]
  wire  _T_4941 = _T_4940 | _T_4814; // @[Mux.scala 27:72]
  wire  _T_4687 = ifu_ic_rw_int_addr_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_17; // @[Reg.scala 27:20]
  wire  _T_4815 = _T_4687 & way_status_out_17; // @[Mux.scala 27:72]
  wire  _T_4942 = _T_4941 | _T_4815; // @[Mux.scala 27:72]
  wire  _T_4688 = ifu_ic_rw_int_addr_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_18; // @[Reg.scala 27:20]
  wire  _T_4816 = _T_4688 & way_status_out_18; // @[Mux.scala 27:72]
  wire  _T_4943 = _T_4942 | _T_4816; // @[Mux.scala 27:72]
  wire  _T_4689 = ifu_ic_rw_int_addr_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_19; // @[Reg.scala 27:20]
  wire  _T_4817 = _T_4689 & way_status_out_19; // @[Mux.scala 27:72]
  wire  _T_4944 = _T_4943 | _T_4817; // @[Mux.scala 27:72]
  wire  _T_4690 = ifu_ic_rw_int_addr_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_20; // @[Reg.scala 27:20]
  wire  _T_4818 = _T_4690 & way_status_out_20; // @[Mux.scala 27:72]
  wire  _T_4945 = _T_4944 | _T_4818; // @[Mux.scala 27:72]
  wire  _T_4691 = ifu_ic_rw_int_addr_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_21; // @[Reg.scala 27:20]
  wire  _T_4819 = _T_4691 & way_status_out_21; // @[Mux.scala 27:72]
  wire  _T_4946 = _T_4945 | _T_4819; // @[Mux.scala 27:72]
  wire  _T_4692 = ifu_ic_rw_int_addr_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_22; // @[Reg.scala 27:20]
  wire  _T_4820 = _T_4692 & way_status_out_22; // @[Mux.scala 27:72]
  wire  _T_4947 = _T_4946 | _T_4820; // @[Mux.scala 27:72]
  wire  _T_4693 = ifu_ic_rw_int_addr_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_23; // @[Reg.scala 27:20]
  wire  _T_4821 = _T_4693 & way_status_out_23; // @[Mux.scala 27:72]
  wire  _T_4948 = _T_4947 | _T_4821; // @[Mux.scala 27:72]
  wire  _T_4694 = ifu_ic_rw_int_addr_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_24; // @[Reg.scala 27:20]
  wire  _T_4822 = _T_4694 & way_status_out_24; // @[Mux.scala 27:72]
  wire  _T_4949 = _T_4948 | _T_4822; // @[Mux.scala 27:72]
  wire  _T_4695 = ifu_ic_rw_int_addr_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_25; // @[Reg.scala 27:20]
  wire  _T_4823 = _T_4695 & way_status_out_25; // @[Mux.scala 27:72]
  wire  _T_4950 = _T_4949 | _T_4823; // @[Mux.scala 27:72]
  wire  _T_4696 = ifu_ic_rw_int_addr_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_26; // @[Reg.scala 27:20]
  wire  _T_4824 = _T_4696 & way_status_out_26; // @[Mux.scala 27:72]
  wire  _T_4951 = _T_4950 | _T_4824; // @[Mux.scala 27:72]
  wire  _T_4697 = ifu_ic_rw_int_addr_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_27; // @[Reg.scala 27:20]
  wire  _T_4825 = _T_4697 & way_status_out_27; // @[Mux.scala 27:72]
  wire  _T_4952 = _T_4951 | _T_4825; // @[Mux.scala 27:72]
  wire  _T_4698 = ifu_ic_rw_int_addr_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_28; // @[Reg.scala 27:20]
  wire  _T_4826 = _T_4698 & way_status_out_28; // @[Mux.scala 27:72]
  wire  _T_4953 = _T_4952 | _T_4826; // @[Mux.scala 27:72]
  wire  _T_4699 = ifu_ic_rw_int_addr_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_29; // @[Reg.scala 27:20]
  wire  _T_4827 = _T_4699 & way_status_out_29; // @[Mux.scala 27:72]
  wire  _T_4954 = _T_4953 | _T_4827; // @[Mux.scala 27:72]
  wire  _T_4700 = ifu_ic_rw_int_addr_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_30; // @[Reg.scala 27:20]
  wire  _T_4828 = _T_4700 & way_status_out_30; // @[Mux.scala 27:72]
  wire  _T_4955 = _T_4954 | _T_4828; // @[Mux.scala 27:72]
  wire  _T_4701 = ifu_ic_rw_int_addr_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_31; // @[Reg.scala 27:20]
  wire  _T_4829 = _T_4701 & way_status_out_31; // @[Mux.scala 27:72]
  wire  _T_4956 = _T_4955 | _T_4829; // @[Mux.scala 27:72]
  wire  _T_4702 = ifu_ic_rw_int_addr_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_32; // @[Reg.scala 27:20]
  wire  _T_4830 = _T_4702 & way_status_out_32; // @[Mux.scala 27:72]
  wire  _T_4957 = _T_4956 | _T_4830; // @[Mux.scala 27:72]
  wire  _T_4703 = ifu_ic_rw_int_addr_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_33; // @[Reg.scala 27:20]
  wire  _T_4831 = _T_4703 & way_status_out_33; // @[Mux.scala 27:72]
  wire  _T_4958 = _T_4957 | _T_4831; // @[Mux.scala 27:72]
  wire  _T_4704 = ifu_ic_rw_int_addr_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_34; // @[Reg.scala 27:20]
  wire  _T_4832 = _T_4704 & way_status_out_34; // @[Mux.scala 27:72]
  wire  _T_4959 = _T_4958 | _T_4832; // @[Mux.scala 27:72]
  wire  _T_4705 = ifu_ic_rw_int_addr_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_35; // @[Reg.scala 27:20]
  wire  _T_4833 = _T_4705 & way_status_out_35; // @[Mux.scala 27:72]
  wire  _T_4960 = _T_4959 | _T_4833; // @[Mux.scala 27:72]
  wire  _T_4706 = ifu_ic_rw_int_addr_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_36; // @[Reg.scala 27:20]
  wire  _T_4834 = _T_4706 & way_status_out_36; // @[Mux.scala 27:72]
  wire  _T_4961 = _T_4960 | _T_4834; // @[Mux.scala 27:72]
  wire  _T_4707 = ifu_ic_rw_int_addr_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_37; // @[Reg.scala 27:20]
  wire  _T_4835 = _T_4707 & way_status_out_37; // @[Mux.scala 27:72]
  wire  _T_4962 = _T_4961 | _T_4835; // @[Mux.scala 27:72]
  wire  _T_4708 = ifu_ic_rw_int_addr_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_38; // @[Reg.scala 27:20]
  wire  _T_4836 = _T_4708 & way_status_out_38; // @[Mux.scala 27:72]
  wire  _T_4963 = _T_4962 | _T_4836; // @[Mux.scala 27:72]
  wire  _T_4709 = ifu_ic_rw_int_addr_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_39; // @[Reg.scala 27:20]
  wire  _T_4837 = _T_4709 & way_status_out_39; // @[Mux.scala 27:72]
  wire  _T_4964 = _T_4963 | _T_4837; // @[Mux.scala 27:72]
  wire  _T_4710 = ifu_ic_rw_int_addr_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_40; // @[Reg.scala 27:20]
  wire  _T_4838 = _T_4710 & way_status_out_40; // @[Mux.scala 27:72]
  wire  _T_4965 = _T_4964 | _T_4838; // @[Mux.scala 27:72]
  wire  _T_4711 = ifu_ic_rw_int_addr_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_41; // @[Reg.scala 27:20]
  wire  _T_4839 = _T_4711 & way_status_out_41; // @[Mux.scala 27:72]
  wire  _T_4966 = _T_4965 | _T_4839; // @[Mux.scala 27:72]
  wire  _T_4712 = ifu_ic_rw_int_addr_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_42; // @[Reg.scala 27:20]
  wire  _T_4840 = _T_4712 & way_status_out_42; // @[Mux.scala 27:72]
  wire  _T_4967 = _T_4966 | _T_4840; // @[Mux.scala 27:72]
  wire  _T_4713 = ifu_ic_rw_int_addr_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_43; // @[Reg.scala 27:20]
  wire  _T_4841 = _T_4713 & way_status_out_43; // @[Mux.scala 27:72]
  wire  _T_4968 = _T_4967 | _T_4841; // @[Mux.scala 27:72]
  wire  _T_4714 = ifu_ic_rw_int_addr_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_44; // @[Reg.scala 27:20]
  wire  _T_4842 = _T_4714 & way_status_out_44; // @[Mux.scala 27:72]
  wire  _T_4969 = _T_4968 | _T_4842; // @[Mux.scala 27:72]
  wire  _T_4715 = ifu_ic_rw_int_addr_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_45; // @[Reg.scala 27:20]
  wire  _T_4843 = _T_4715 & way_status_out_45; // @[Mux.scala 27:72]
  wire  _T_4970 = _T_4969 | _T_4843; // @[Mux.scala 27:72]
  wire  _T_4716 = ifu_ic_rw_int_addr_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_46; // @[Reg.scala 27:20]
  wire  _T_4844 = _T_4716 & way_status_out_46; // @[Mux.scala 27:72]
  wire  _T_4971 = _T_4970 | _T_4844; // @[Mux.scala 27:72]
  wire  _T_4717 = ifu_ic_rw_int_addr_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_47; // @[Reg.scala 27:20]
  wire  _T_4845 = _T_4717 & way_status_out_47; // @[Mux.scala 27:72]
  wire  _T_4972 = _T_4971 | _T_4845; // @[Mux.scala 27:72]
  wire  _T_4718 = ifu_ic_rw_int_addr_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_48; // @[Reg.scala 27:20]
  wire  _T_4846 = _T_4718 & way_status_out_48; // @[Mux.scala 27:72]
  wire  _T_4973 = _T_4972 | _T_4846; // @[Mux.scala 27:72]
  wire  _T_4719 = ifu_ic_rw_int_addr_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_49; // @[Reg.scala 27:20]
  wire  _T_4847 = _T_4719 & way_status_out_49; // @[Mux.scala 27:72]
  wire  _T_4974 = _T_4973 | _T_4847; // @[Mux.scala 27:72]
  wire  _T_4720 = ifu_ic_rw_int_addr_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_50; // @[Reg.scala 27:20]
  wire  _T_4848 = _T_4720 & way_status_out_50; // @[Mux.scala 27:72]
  wire  _T_4975 = _T_4974 | _T_4848; // @[Mux.scala 27:72]
  wire  _T_4721 = ifu_ic_rw_int_addr_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_51; // @[Reg.scala 27:20]
  wire  _T_4849 = _T_4721 & way_status_out_51; // @[Mux.scala 27:72]
  wire  _T_4976 = _T_4975 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4722 = ifu_ic_rw_int_addr_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_52; // @[Reg.scala 27:20]
  wire  _T_4850 = _T_4722 & way_status_out_52; // @[Mux.scala 27:72]
  wire  _T_4977 = _T_4976 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4723 = ifu_ic_rw_int_addr_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_53; // @[Reg.scala 27:20]
  wire  _T_4851 = _T_4723 & way_status_out_53; // @[Mux.scala 27:72]
  wire  _T_4978 = _T_4977 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_4724 = ifu_ic_rw_int_addr_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_54; // @[Reg.scala 27:20]
  wire  _T_4852 = _T_4724 & way_status_out_54; // @[Mux.scala 27:72]
  wire  _T_4979 = _T_4978 | _T_4852; // @[Mux.scala 27:72]
  wire  _T_4725 = ifu_ic_rw_int_addr_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_55; // @[Reg.scala 27:20]
  wire  _T_4853 = _T_4725 & way_status_out_55; // @[Mux.scala 27:72]
  wire  _T_4980 = _T_4979 | _T_4853; // @[Mux.scala 27:72]
  wire  _T_4726 = ifu_ic_rw_int_addr_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_56; // @[Reg.scala 27:20]
  wire  _T_4854 = _T_4726 & way_status_out_56; // @[Mux.scala 27:72]
  wire  _T_4981 = _T_4980 | _T_4854; // @[Mux.scala 27:72]
  wire  _T_4727 = ifu_ic_rw_int_addr_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_57; // @[Reg.scala 27:20]
  wire  _T_4855 = _T_4727 & way_status_out_57; // @[Mux.scala 27:72]
  wire  _T_4982 = _T_4981 | _T_4855; // @[Mux.scala 27:72]
  wire  _T_4728 = ifu_ic_rw_int_addr_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_58; // @[Reg.scala 27:20]
  wire  _T_4856 = _T_4728 & way_status_out_58; // @[Mux.scala 27:72]
  wire  _T_4983 = _T_4982 | _T_4856; // @[Mux.scala 27:72]
  wire  _T_4729 = ifu_ic_rw_int_addr_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_59; // @[Reg.scala 27:20]
  wire  _T_4857 = _T_4729 & way_status_out_59; // @[Mux.scala 27:72]
  wire  _T_4984 = _T_4983 | _T_4857; // @[Mux.scala 27:72]
  wire  _T_4730 = ifu_ic_rw_int_addr_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_60; // @[Reg.scala 27:20]
  wire  _T_4858 = _T_4730 & way_status_out_60; // @[Mux.scala 27:72]
  wire  _T_4985 = _T_4984 | _T_4858; // @[Mux.scala 27:72]
  wire  _T_4731 = ifu_ic_rw_int_addr_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_61; // @[Reg.scala 27:20]
  wire  _T_4859 = _T_4731 & way_status_out_61; // @[Mux.scala 27:72]
  wire  _T_4986 = _T_4985 | _T_4859; // @[Mux.scala 27:72]
  wire  _T_4732 = ifu_ic_rw_int_addr_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_62; // @[Reg.scala 27:20]
  wire  _T_4860 = _T_4732 & way_status_out_62; // @[Mux.scala 27:72]
  wire  _T_4987 = _T_4986 | _T_4860; // @[Mux.scala 27:72]
  wire  _T_4733 = ifu_ic_rw_int_addr_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_63; // @[Reg.scala 27:20]
  wire  _T_4861 = _T_4733 & way_status_out_63; // @[Mux.scala 27:72]
  wire  _T_4988 = _T_4987 | _T_4861; // @[Mux.scala 27:72]
  wire  _T_4734 = ifu_ic_rw_int_addr_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_64; // @[Reg.scala 27:20]
  wire  _T_4862 = _T_4734 & way_status_out_64; // @[Mux.scala 27:72]
  wire  _T_4989 = _T_4988 | _T_4862; // @[Mux.scala 27:72]
  wire  _T_4735 = ifu_ic_rw_int_addr_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_65; // @[Reg.scala 27:20]
  wire  _T_4863 = _T_4735 & way_status_out_65; // @[Mux.scala 27:72]
  wire  _T_4990 = _T_4989 | _T_4863; // @[Mux.scala 27:72]
  wire  _T_4736 = ifu_ic_rw_int_addr_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_66; // @[Reg.scala 27:20]
  wire  _T_4864 = _T_4736 & way_status_out_66; // @[Mux.scala 27:72]
  wire  _T_4991 = _T_4990 | _T_4864; // @[Mux.scala 27:72]
  wire  _T_4737 = ifu_ic_rw_int_addr_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_67; // @[Reg.scala 27:20]
  wire  _T_4865 = _T_4737 & way_status_out_67; // @[Mux.scala 27:72]
  wire  _T_4992 = _T_4991 | _T_4865; // @[Mux.scala 27:72]
  wire  _T_4738 = ifu_ic_rw_int_addr_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_68; // @[Reg.scala 27:20]
  wire  _T_4866 = _T_4738 & way_status_out_68; // @[Mux.scala 27:72]
  wire  _T_4993 = _T_4992 | _T_4866; // @[Mux.scala 27:72]
  wire  _T_4739 = ifu_ic_rw_int_addr_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_69; // @[Reg.scala 27:20]
  wire  _T_4867 = _T_4739 & way_status_out_69; // @[Mux.scala 27:72]
  wire  _T_4994 = _T_4993 | _T_4867; // @[Mux.scala 27:72]
  wire  _T_4740 = ifu_ic_rw_int_addr_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_70; // @[Reg.scala 27:20]
  wire  _T_4868 = _T_4740 & way_status_out_70; // @[Mux.scala 27:72]
  wire  _T_4995 = _T_4994 | _T_4868; // @[Mux.scala 27:72]
  wire  _T_4741 = ifu_ic_rw_int_addr_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_71; // @[Reg.scala 27:20]
  wire  _T_4869 = _T_4741 & way_status_out_71; // @[Mux.scala 27:72]
  wire  _T_4996 = _T_4995 | _T_4869; // @[Mux.scala 27:72]
  wire  _T_4742 = ifu_ic_rw_int_addr_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_72; // @[Reg.scala 27:20]
  wire  _T_4870 = _T_4742 & way_status_out_72; // @[Mux.scala 27:72]
  wire  _T_4997 = _T_4996 | _T_4870; // @[Mux.scala 27:72]
  wire  _T_4743 = ifu_ic_rw_int_addr_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_73; // @[Reg.scala 27:20]
  wire  _T_4871 = _T_4743 & way_status_out_73; // @[Mux.scala 27:72]
  wire  _T_4998 = _T_4997 | _T_4871; // @[Mux.scala 27:72]
  wire  _T_4744 = ifu_ic_rw_int_addr_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_74; // @[Reg.scala 27:20]
  wire  _T_4872 = _T_4744 & way_status_out_74; // @[Mux.scala 27:72]
  wire  _T_4999 = _T_4998 | _T_4872; // @[Mux.scala 27:72]
  wire  _T_4745 = ifu_ic_rw_int_addr_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_75; // @[Reg.scala 27:20]
  wire  _T_4873 = _T_4745 & way_status_out_75; // @[Mux.scala 27:72]
  wire  _T_5000 = _T_4999 | _T_4873; // @[Mux.scala 27:72]
  wire  _T_4746 = ifu_ic_rw_int_addr_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_76; // @[Reg.scala 27:20]
  wire  _T_4874 = _T_4746 & way_status_out_76; // @[Mux.scala 27:72]
  wire  _T_5001 = _T_5000 | _T_4874; // @[Mux.scala 27:72]
  wire  _T_4747 = ifu_ic_rw_int_addr_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_77; // @[Reg.scala 27:20]
  wire  _T_4875 = _T_4747 & way_status_out_77; // @[Mux.scala 27:72]
  wire  _T_5002 = _T_5001 | _T_4875; // @[Mux.scala 27:72]
  wire  _T_4748 = ifu_ic_rw_int_addr_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_78; // @[Reg.scala 27:20]
  wire  _T_4876 = _T_4748 & way_status_out_78; // @[Mux.scala 27:72]
  wire  _T_5003 = _T_5002 | _T_4876; // @[Mux.scala 27:72]
  wire  _T_4749 = ifu_ic_rw_int_addr_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_79; // @[Reg.scala 27:20]
  wire  _T_4877 = _T_4749 & way_status_out_79; // @[Mux.scala 27:72]
  wire  _T_5004 = _T_5003 | _T_4877; // @[Mux.scala 27:72]
  wire  _T_4750 = ifu_ic_rw_int_addr_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_80; // @[Reg.scala 27:20]
  wire  _T_4878 = _T_4750 & way_status_out_80; // @[Mux.scala 27:72]
  wire  _T_5005 = _T_5004 | _T_4878; // @[Mux.scala 27:72]
  wire  _T_4751 = ifu_ic_rw_int_addr_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_81; // @[Reg.scala 27:20]
  wire  _T_4879 = _T_4751 & way_status_out_81; // @[Mux.scala 27:72]
  wire  _T_5006 = _T_5005 | _T_4879; // @[Mux.scala 27:72]
  wire  _T_4752 = ifu_ic_rw_int_addr_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_82; // @[Reg.scala 27:20]
  wire  _T_4880 = _T_4752 & way_status_out_82; // @[Mux.scala 27:72]
  wire  _T_5007 = _T_5006 | _T_4880; // @[Mux.scala 27:72]
  wire  _T_4753 = ifu_ic_rw_int_addr_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_83; // @[Reg.scala 27:20]
  wire  _T_4881 = _T_4753 & way_status_out_83; // @[Mux.scala 27:72]
  wire  _T_5008 = _T_5007 | _T_4881; // @[Mux.scala 27:72]
  wire  _T_4754 = ifu_ic_rw_int_addr_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_84; // @[Reg.scala 27:20]
  wire  _T_4882 = _T_4754 & way_status_out_84; // @[Mux.scala 27:72]
  wire  _T_5009 = _T_5008 | _T_4882; // @[Mux.scala 27:72]
  wire  _T_4755 = ifu_ic_rw_int_addr_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_85; // @[Reg.scala 27:20]
  wire  _T_4883 = _T_4755 & way_status_out_85; // @[Mux.scala 27:72]
  wire  _T_5010 = _T_5009 | _T_4883; // @[Mux.scala 27:72]
  wire  _T_4756 = ifu_ic_rw_int_addr_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_86; // @[Reg.scala 27:20]
  wire  _T_4884 = _T_4756 & way_status_out_86; // @[Mux.scala 27:72]
  wire  _T_5011 = _T_5010 | _T_4884; // @[Mux.scala 27:72]
  wire  _T_4757 = ifu_ic_rw_int_addr_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_87; // @[Reg.scala 27:20]
  wire  _T_4885 = _T_4757 & way_status_out_87; // @[Mux.scala 27:72]
  wire  _T_5012 = _T_5011 | _T_4885; // @[Mux.scala 27:72]
  wire  _T_4758 = ifu_ic_rw_int_addr_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_88; // @[Reg.scala 27:20]
  wire  _T_4886 = _T_4758 & way_status_out_88; // @[Mux.scala 27:72]
  wire  _T_5013 = _T_5012 | _T_4886; // @[Mux.scala 27:72]
  wire  _T_4759 = ifu_ic_rw_int_addr_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_89; // @[Reg.scala 27:20]
  wire  _T_4887 = _T_4759 & way_status_out_89; // @[Mux.scala 27:72]
  wire  _T_5014 = _T_5013 | _T_4887; // @[Mux.scala 27:72]
  wire  _T_4760 = ifu_ic_rw_int_addr_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_90; // @[Reg.scala 27:20]
  wire  _T_4888 = _T_4760 & way_status_out_90; // @[Mux.scala 27:72]
  wire  _T_5015 = _T_5014 | _T_4888; // @[Mux.scala 27:72]
  wire  _T_4761 = ifu_ic_rw_int_addr_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_91; // @[Reg.scala 27:20]
  wire  _T_4889 = _T_4761 & way_status_out_91; // @[Mux.scala 27:72]
  wire  _T_5016 = _T_5015 | _T_4889; // @[Mux.scala 27:72]
  wire  _T_4762 = ifu_ic_rw_int_addr_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_92; // @[Reg.scala 27:20]
  wire  _T_4890 = _T_4762 & way_status_out_92; // @[Mux.scala 27:72]
  wire  _T_5017 = _T_5016 | _T_4890; // @[Mux.scala 27:72]
  wire  _T_4763 = ifu_ic_rw_int_addr_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_93; // @[Reg.scala 27:20]
  wire  _T_4891 = _T_4763 & way_status_out_93; // @[Mux.scala 27:72]
  wire  _T_5018 = _T_5017 | _T_4891; // @[Mux.scala 27:72]
  wire  _T_4764 = ifu_ic_rw_int_addr_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_94; // @[Reg.scala 27:20]
  wire  _T_4892 = _T_4764 & way_status_out_94; // @[Mux.scala 27:72]
  wire  _T_5019 = _T_5018 | _T_4892; // @[Mux.scala 27:72]
  wire  _T_4765 = ifu_ic_rw_int_addr_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_95; // @[Reg.scala 27:20]
  wire  _T_4893 = _T_4765 & way_status_out_95; // @[Mux.scala 27:72]
  wire  _T_5020 = _T_5019 | _T_4893; // @[Mux.scala 27:72]
  wire  _T_4766 = ifu_ic_rw_int_addr_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_96; // @[Reg.scala 27:20]
  wire  _T_4894 = _T_4766 & way_status_out_96; // @[Mux.scala 27:72]
  wire  _T_5021 = _T_5020 | _T_4894; // @[Mux.scala 27:72]
  wire  _T_4767 = ifu_ic_rw_int_addr_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_97; // @[Reg.scala 27:20]
  wire  _T_4895 = _T_4767 & way_status_out_97; // @[Mux.scala 27:72]
  wire  _T_5022 = _T_5021 | _T_4895; // @[Mux.scala 27:72]
  wire  _T_4768 = ifu_ic_rw_int_addr_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_98; // @[Reg.scala 27:20]
  wire  _T_4896 = _T_4768 & way_status_out_98; // @[Mux.scala 27:72]
  wire  _T_5023 = _T_5022 | _T_4896; // @[Mux.scala 27:72]
  wire  _T_4769 = ifu_ic_rw_int_addr_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_99; // @[Reg.scala 27:20]
  wire  _T_4897 = _T_4769 & way_status_out_99; // @[Mux.scala 27:72]
  wire  _T_5024 = _T_5023 | _T_4897; // @[Mux.scala 27:72]
  wire  _T_4770 = ifu_ic_rw_int_addr_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_100; // @[Reg.scala 27:20]
  wire  _T_4898 = _T_4770 & way_status_out_100; // @[Mux.scala 27:72]
  wire  _T_5025 = _T_5024 | _T_4898; // @[Mux.scala 27:72]
  wire  _T_4771 = ifu_ic_rw_int_addr_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_101; // @[Reg.scala 27:20]
  wire  _T_4899 = _T_4771 & way_status_out_101; // @[Mux.scala 27:72]
  wire  _T_5026 = _T_5025 | _T_4899; // @[Mux.scala 27:72]
  wire  _T_4772 = ifu_ic_rw_int_addr_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_102; // @[Reg.scala 27:20]
  wire  _T_4900 = _T_4772 & way_status_out_102; // @[Mux.scala 27:72]
  wire  _T_5027 = _T_5026 | _T_4900; // @[Mux.scala 27:72]
  wire  _T_4773 = ifu_ic_rw_int_addr_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_103; // @[Reg.scala 27:20]
  wire  _T_4901 = _T_4773 & way_status_out_103; // @[Mux.scala 27:72]
  wire  _T_5028 = _T_5027 | _T_4901; // @[Mux.scala 27:72]
  wire  _T_4774 = ifu_ic_rw_int_addr_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_104; // @[Reg.scala 27:20]
  wire  _T_4902 = _T_4774 & way_status_out_104; // @[Mux.scala 27:72]
  wire  _T_5029 = _T_5028 | _T_4902; // @[Mux.scala 27:72]
  wire  _T_4775 = ifu_ic_rw_int_addr_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_105; // @[Reg.scala 27:20]
  wire  _T_4903 = _T_4775 & way_status_out_105; // @[Mux.scala 27:72]
  wire  _T_5030 = _T_5029 | _T_4903; // @[Mux.scala 27:72]
  wire  _T_4776 = ifu_ic_rw_int_addr_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_106; // @[Reg.scala 27:20]
  wire  _T_4904 = _T_4776 & way_status_out_106; // @[Mux.scala 27:72]
  wire  _T_5031 = _T_5030 | _T_4904; // @[Mux.scala 27:72]
  wire  _T_4777 = ifu_ic_rw_int_addr_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_107; // @[Reg.scala 27:20]
  wire  _T_4905 = _T_4777 & way_status_out_107; // @[Mux.scala 27:72]
  wire  _T_5032 = _T_5031 | _T_4905; // @[Mux.scala 27:72]
  wire  _T_4778 = ifu_ic_rw_int_addr_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_108; // @[Reg.scala 27:20]
  wire  _T_4906 = _T_4778 & way_status_out_108; // @[Mux.scala 27:72]
  wire  _T_5033 = _T_5032 | _T_4906; // @[Mux.scala 27:72]
  wire  _T_4779 = ifu_ic_rw_int_addr_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_109; // @[Reg.scala 27:20]
  wire  _T_4907 = _T_4779 & way_status_out_109; // @[Mux.scala 27:72]
  wire  _T_5034 = _T_5033 | _T_4907; // @[Mux.scala 27:72]
  wire  _T_4780 = ifu_ic_rw_int_addr_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_110; // @[Reg.scala 27:20]
  wire  _T_4908 = _T_4780 & way_status_out_110; // @[Mux.scala 27:72]
  wire  _T_5035 = _T_5034 | _T_4908; // @[Mux.scala 27:72]
  wire  _T_4781 = ifu_ic_rw_int_addr_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_111; // @[Reg.scala 27:20]
  wire  _T_4909 = _T_4781 & way_status_out_111; // @[Mux.scala 27:72]
  wire  _T_5036 = _T_5035 | _T_4909; // @[Mux.scala 27:72]
  wire  _T_4782 = ifu_ic_rw_int_addr_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_112; // @[Reg.scala 27:20]
  wire  _T_4910 = _T_4782 & way_status_out_112; // @[Mux.scala 27:72]
  wire  _T_5037 = _T_5036 | _T_4910; // @[Mux.scala 27:72]
  wire  _T_4783 = ifu_ic_rw_int_addr_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_113; // @[Reg.scala 27:20]
  wire  _T_4911 = _T_4783 & way_status_out_113; // @[Mux.scala 27:72]
  wire  _T_5038 = _T_5037 | _T_4911; // @[Mux.scala 27:72]
  wire  _T_4784 = ifu_ic_rw_int_addr_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_114; // @[Reg.scala 27:20]
  wire  _T_4912 = _T_4784 & way_status_out_114; // @[Mux.scala 27:72]
  wire  _T_5039 = _T_5038 | _T_4912; // @[Mux.scala 27:72]
  wire  _T_4785 = ifu_ic_rw_int_addr_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_115; // @[Reg.scala 27:20]
  wire  _T_4913 = _T_4785 & way_status_out_115; // @[Mux.scala 27:72]
  wire  _T_5040 = _T_5039 | _T_4913; // @[Mux.scala 27:72]
  wire  _T_4786 = ifu_ic_rw_int_addr_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_116; // @[Reg.scala 27:20]
  wire  _T_4914 = _T_4786 & way_status_out_116; // @[Mux.scala 27:72]
  wire  _T_5041 = _T_5040 | _T_4914; // @[Mux.scala 27:72]
  wire  _T_4787 = ifu_ic_rw_int_addr_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_117; // @[Reg.scala 27:20]
  wire  _T_4915 = _T_4787 & way_status_out_117; // @[Mux.scala 27:72]
  wire  _T_5042 = _T_5041 | _T_4915; // @[Mux.scala 27:72]
  wire  _T_4788 = ifu_ic_rw_int_addr_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_118; // @[Reg.scala 27:20]
  wire  _T_4916 = _T_4788 & way_status_out_118; // @[Mux.scala 27:72]
  wire  _T_5043 = _T_5042 | _T_4916; // @[Mux.scala 27:72]
  wire  _T_4789 = ifu_ic_rw_int_addr_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_119; // @[Reg.scala 27:20]
  wire  _T_4917 = _T_4789 & way_status_out_119; // @[Mux.scala 27:72]
  wire  _T_5044 = _T_5043 | _T_4917; // @[Mux.scala 27:72]
  wire  _T_4790 = ifu_ic_rw_int_addr_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_120; // @[Reg.scala 27:20]
  wire  _T_4918 = _T_4790 & way_status_out_120; // @[Mux.scala 27:72]
  wire  _T_5045 = _T_5044 | _T_4918; // @[Mux.scala 27:72]
  wire  _T_4791 = ifu_ic_rw_int_addr_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_121; // @[Reg.scala 27:20]
  wire  _T_4919 = _T_4791 & way_status_out_121; // @[Mux.scala 27:72]
  wire  _T_5046 = _T_5045 | _T_4919; // @[Mux.scala 27:72]
  wire  _T_4792 = ifu_ic_rw_int_addr_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_122; // @[Reg.scala 27:20]
  wire  _T_4920 = _T_4792 & way_status_out_122; // @[Mux.scala 27:72]
  wire  _T_5047 = _T_5046 | _T_4920; // @[Mux.scala 27:72]
  wire  _T_4793 = ifu_ic_rw_int_addr_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_123; // @[Reg.scala 27:20]
  wire  _T_4921 = _T_4793 & way_status_out_123; // @[Mux.scala 27:72]
  wire  _T_5048 = _T_5047 | _T_4921; // @[Mux.scala 27:72]
  wire  _T_4794 = ifu_ic_rw_int_addr_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_124; // @[Reg.scala 27:20]
  wire  _T_4922 = _T_4794 & way_status_out_124; // @[Mux.scala 27:72]
  wire  _T_5049 = _T_5048 | _T_4922; // @[Mux.scala 27:72]
  wire  _T_4795 = ifu_ic_rw_int_addr_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_125; // @[Reg.scala 27:20]
  wire  _T_4923 = _T_4795 & way_status_out_125; // @[Mux.scala 27:72]
  wire  _T_5050 = _T_5049 | _T_4923; // @[Mux.scala 27:72]
  wire  _T_4796 = ifu_ic_rw_int_addr_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_126; // @[Reg.scala 27:20]
  wire  _T_4924 = _T_4796 & way_status_out_126; // @[Mux.scala 27:72]
  wire  _T_5051 = _T_5050 | _T_4924; // @[Mux.scala 27:72]
  wire  _T_4797 = ifu_ic_rw_int_addr_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 738:80]
  reg  way_status_out_127; // @[Reg.scala 27:20]
  wire  _T_4925 = _T_4797 & way_status_out_127; // @[Mux.scala 27:72]
  wire  way_status = _T_5051 | _T_4925; // @[Mux.scala 27:72]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 263:96]
  wire [1:0] _T_197 = _T_195 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_198 = _T_197 & io_ic_tag_valid; // @[el2_ifu_mem_ctl.scala 263:113]
  reg [1:0] tagv_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 269:58]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 265:67]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 267:54]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[el2_ifu_mem_ctl.scala 588:46]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 272:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 277:59]
  wire  _T_214 = _T_212 | _T_2267; // @[el2_ifu_mem_ctl.scala 277:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 277:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 283:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 283:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 283:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 283:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 290:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 290:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 290:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 291:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 291:32]
  wire  _T_274 = imb_ff[11:5] == imb_scnd_ff[11:5]; // @[el2_ifu_mem_ctl.scala 294:79]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 294:135]
  reg [1:0] ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 586:51]
  wire  _T_2692 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 631:48]
  wire  _T_2693 = _T_2692 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 631:52]
  wire  bus_ifu_wr_data_error_ff = _T_2693 & miss_pending; // @[el2_ifu_mem_ctl.scala 631:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 368:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 367:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 294:153]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 294:151]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 297:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 297:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 298:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 318:59]
  wire  _T_9755 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 794:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 319:53]
  wire  _T_9757 = _T_9755 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 794:51]
  wire  _T_9759 = _T_9757 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 794:67]
  wire  _T_9761 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 794:86]
  wire  replace_way_mb_any_0 = _T_9759 | _T_9761; // @[el2_ifu_mem_ctl.scala 794:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9764 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 795:50]
  wire  _T_9766 = _T_9764 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 795:66]
  wire  _T_9768 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 795:85]
  wire  _T_9770 = _T_9768 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 795:100]
  wire  replace_way_mb_any_1 = _T_9766 | _T_9770; // @[el2_ifu_mem_ctl.scala 795:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 302:110]
  wire [1:0] _T_290 = tagv_mb_scnd_ff | _T_289; // @[el2_ifu_mem_ctl.scala 302:62]
  wire [1:0] _T_295 = io_ic_tag_valid & _T_197; // @[el2_ifu_mem_ctl.scala 303:56]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 306:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 306:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 307:48]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 306:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 306:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 308:62]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 317:48]
  wire  _T_309 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 316:57]
  wire  _T_315 = _T_2282 & flush_final_f; // @[el2_ifu_mem_ctl.scala 321:87]
  wire  _T_316 = ~_T_315; // @[el2_ifu_mem_ctl.scala 321:55]
  wire  _T_317 = io_ifc_fetch_req_bf & _T_316; // @[el2_ifu_mem_ctl.scala 321:53]
  wire  _T_2274 = ~_T_2269; // @[el2_ifu_mem_ctl.scala 466:46]
  wire  _T_2275 = _T_2267 & _T_2274; // @[el2_ifu_mem_ctl.scala 466:44]
  wire  stream_miss_f = _T_2275 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 466:84]
  wire  _T_318 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 321:106]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 327:68]
  reg [2:0] bus_rd_addr_count; // @[el2_ifu_mem_ctl.scala 613:55]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_325 = _T_239 | _T_2267; // @[el2_ifu_mem_ctl.scala 329:55]
  wire  _T_328 = _T_325 & _T_56; // @[el2_ifu_mem_ctl.scala 329:82]
  wire  _T_2288 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 471:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2288}; // @[Cat.scala 29:58]
  wire  _T_2289 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 472:81]
  wire  _T_2313 = _T_2289 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2292 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 472:81]
  wire  _T_2314 = _T_2292 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2321 = _T_2313 | _T_2314; // @[Mux.scala 27:72]
  wire  _T_2295 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 472:81]
  wire  _T_2315 = _T_2295 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2322 = _T_2321 | _T_2315; // @[Mux.scala 27:72]
  wire  _T_2298 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 472:81]
  wire  _T_2316 = _T_2298 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2323 = _T_2322 | _T_2316; // @[Mux.scala 27:72]
  wire  _T_2301 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 472:81]
  wire  _T_2317 = _T_2301 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2324 = _T_2323 | _T_2317; // @[Mux.scala 27:72]
  wire  _T_2304 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 472:81]
  wire  _T_2318 = _T_2304 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2325 = _T_2324 | _T_2318; // @[Mux.scala 27:72]
  wire  _T_2307 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 472:81]
  wire  _T_2319 = _T_2307 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2326 = _T_2325 | _T_2319; // @[Mux.scala 27:72]
  wire  _T_2310 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 472:81]
  wire  _T_2320 = _T_2310 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2326 | _T_2320; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 473:46]
  wire  _T_332 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 333:35]
  wire  _T_334 = _T_332 & _T_17; // @[el2_ifu_mem_ctl.scala 333:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 628:61]
  wire  _T_2686 = ic_act_miss_f_delayed & _T_2283; // @[el2_ifu_mem_ctl.scala 629:53]
  wire  reset_tag_valid_for_miss = _T_2686 & _T_17; // @[el2_ifu_mem_ctl.scala 629:84]
  wire  sel_mb_addr = _T_334 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 333:79]
  wire [30:0] _T_338 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_339 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 335:37]
  wire [30:0] _T_340 = sel_mb_addr ? _T_338 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_341 = _T_339 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_340 | _T_341; // @[Mux.scala 27:72]
  wire  _T_346 = _T_334 & last_beat; // @[el2_ifu_mem_ctl.scala 337:84]
  wire  _T_2680 = ~_T_2692; // @[el2_ifu_mem_ctl.scala 626:84]
  wire  _T_2681 = _T_100 & _T_2680; // @[el2_ifu_mem_ctl.scala 626:82]
  wire  bus_ifu_wr_en_ff_q = _T_2681 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 626:108]
  wire  sel_mb_status_addr = _T_346 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 337:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_338 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 338:31]
  reg [63:0] ifu_bus_rdata_ff; // @[el2_ifu_mem_ctl.scala 587:48]
  wire [6:0] _T_569 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 416:13]
  wire  _T_570 = ^_T_569; // @[el2_lib.scala 416:20]
  wire [6:0] _T_576 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_583 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 416:30]
  wire [14:0] _T_584 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_576}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_591 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 416:30]
  wire [30:0] _T_600 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_591,_T_584}; // @[el2_lib.scala 416:30]
  wire  _T_601 = ^_T_600; // @[el2_lib.scala 416:37]
  wire [6:0] _T_607 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 416:47]
  wire [14:0] _T_615 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_607}; // @[el2_lib.scala 416:47]
  wire [30:0] _T_631 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_591,_T_615}; // @[el2_lib.scala 416:47]
  wire  _T_632 = ^_T_631; // @[el2_lib.scala 416:54]
  wire [6:0] _T_638 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 416:64]
  wire [14:0] _T_646 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_638}; // @[el2_lib.scala 416:64]
  wire [30:0] _T_662 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_583,_T_646}; // @[el2_lib.scala 416:64]
  wire  _T_663 = ^_T_662; // @[el2_lib.scala 416:71]
  wire [7:0] _T_670 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 416:81]
  wire [16:0] _T_679 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_670}; // @[el2_lib.scala 416:81]
  wire [8:0] _T_687 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 416:81]
  wire [17:0] _T_696 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_687}; // @[el2_lib.scala 416:81]
  wire [34:0] _T_697 = {_T_696,_T_679}; // @[el2_lib.scala 416:81]
  wire  _T_698 = ^_T_697; // @[el2_lib.scala 416:88]
  wire [7:0] _T_705 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 416:98]
  wire [16:0] _T_714 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_705}; // @[el2_lib.scala 416:98]
  wire [8:0] _T_722 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 416:98]
  wire [17:0] _T_731 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_722}; // @[el2_lib.scala 416:98]
  wire [34:0] _T_732 = {_T_731,_T_714}; // @[el2_lib.scala 416:98]
  wire  _T_733 = ^_T_732; // @[el2_lib.scala 416:105]
  wire [7:0] _T_740 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 416:115]
  wire [16:0] _T_749 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_740}; // @[el2_lib.scala 416:115]
  wire [8:0] _T_757 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 416:115]
  wire [17:0] _T_766 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_757}; // @[el2_lib.scala 416:115]
  wire [34:0] _T_767 = {_T_766,_T_749}; // @[el2_lib.scala 416:115]
  wire  _T_768 = ^_T_767; // @[el2_lib.scala 416:122]
  wire [3:0] _T_2329 = {ifu_bus_rid_ff[2:1],_T_2288,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2330 = _T_2329 == 4'h0; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_0; // @[el2_ifu_mem_ctl.scala 408:65]
  wire [31:0] _T_2377 = _T_2330 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2333 = _T_2329 == 4'h1; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_1; // @[el2_ifu_mem_ctl.scala 409:67]
  wire [31:0] _T_2378 = _T_2333 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2393 = _T_2377 | _T_2378; // @[Mux.scala 27:72]
  wire  _T_2336 = _T_2329 == 4'h2; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_2; // @[el2_ifu_mem_ctl.scala 408:65]
  wire [31:0] _T_2379 = _T_2336 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2394 = _T_2393 | _T_2379; // @[Mux.scala 27:72]
  wire  _T_2339 = _T_2329 == 4'h3; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_3; // @[el2_ifu_mem_ctl.scala 409:67]
  wire [31:0] _T_2380 = _T_2339 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2395 = _T_2394 | _T_2380; // @[Mux.scala 27:72]
  wire  _T_2342 = _T_2329 == 4'h4; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_4; // @[el2_ifu_mem_ctl.scala 408:65]
  wire [31:0] _T_2381 = _T_2342 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2396 = _T_2395 | _T_2381; // @[Mux.scala 27:72]
  wire  _T_2345 = _T_2329 == 4'h5; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_5; // @[el2_ifu_mem_ctl.scala 409:67]
  wire [31:0] _T_2382 = _T_2345 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2397 = _T_2396 | _T_2382; // @[Mux.scala 27:72]
  wire  _T_2348 = _T_2329 == 4'h6; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_6; // @[el2_ifu_mem_ctl.scala 408:65]
  wire [31:0] _T_2383 = _T_2348 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2398 = _T_2397 | _T_2383; // @[Mux.scala 27:72]
  wire  _T_2351 = _T_2329 == 4'h7; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_7; // @[el2_ifu_mem_ctl.scala 409:67]
  wire [31:0] _T_2384 = _T_2351 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2399 = _T_2398 | _T_2384; // @[Mux.scala 27:72]
  wire  _T_2354 = _T_2329 == 4'h8; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_8; // @[el2_ifu_mem_ctl.scala 408:65]
  wire [31:0] _T_2385 = _T_2354 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2400 = _T_2399 | _T_2385; // @[Mux.scala 27:72]
  wire  _T_2357 = _T_2329 == 4'h9; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_9; // @[el2_ifu_mem_ctl.scala 409:67]
  wire [31:0] _T_2386 = _T_2357 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2401 = _T_2400 | _T_2386; // @[Mux.scala 27:72]
  wire  _T_2360 = _T_2329 == 4'ha; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_10; // @[el2_ifu_mem_ctl.scala 408:65]
  wire [31:0] _T_2387 = _T_2360 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2402 = _T_2401 | _T_2387; // @[Mux.scala 27:72]
  wire  _T_2363 = _T_2329 == 4'hb; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_11; // @[el2_ifu_mem_ctl.scala 409:67]
  wire [31:0] _T_2388 = _T_2363 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2403 = _T_2402 | _T_2388; // @[Mux.scala 27:72]
  wire  _T_2366 = _T_2329 == 4'hc; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_12; // @[el2_ifu_mem_ctl.scala 408:65]
  wire [31:0] _T_2389 = _T_2366 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2404 = _T_2403 | _T_2389; // @[Mux.scala 27:72]
  wire  _T_2369 = _T_2329 == 4'hd; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_13; // @[el2_ifu_mem_ctl.scala 409:67]
  wire [31:0] _T_2390 = _T_2369 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2405 = _T_2404 | _T_2390; // @[Mux.scala 27:72]
  wire  _T_2372 = _T_2329 == 4'he; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_14; // @[el2_ifu_mem_ctl.scala 408:65]
  wire [31:0] _T_2391 = _T_2372 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2406 = _T_2405 | _T_2391; // @[Mux.scala 27:72]
  wire  _T_2375 = _T_2329 == 4'hf; // @[el2_ifu_mem_ctl.scala 474:89]
  reg [31:0] ic_miss_buff_data_15; // @[el2_ifu_mem_ctl.scala 409:67]
  wire [31:0] _T_2392 = _T_2375 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2407 = _T_2406 | _T_2392; // @[Mux.scala 27:72]
  wire [3:0] _T_2409 = {ifu_bus_rid_ff[2:1],_T_2288,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2410 = _T_2409 == 4'h0; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2457 = _T_2410 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2413 = _T_2409 == 4'h1; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2458 = _T_2413 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2473 = _T_2457 | _T_2458; // @[Mux.scala 27:72]
  wire  _T_2416 = _T_2409 == 4'h2; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2459 = _T_2416 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2474 = _T_2473 | _T_2459; // @[Mux.scala 27:72]
  wire  _T_2419 = _T_2409 == 4'h3; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2460 = _T_2419 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2475 = _T_2474 | _T_2460; // @[Mux.scala 27:72]
  wire  _T_2422 = _T_2409 == 4'h4; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2461 = _T_2422 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2476 = _T_2475 | _T_2461; // @[Mux.scala 27:72]
  wire  _T_2425 = _T_2409 == 4'h5; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2462 = _T_2425 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2477 = _T_2476 | _T_2462; // @[Mux.scala 27:72]
  wire  _T_2428 = _T_2409 == 4'h6; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2463 = _T_2428 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2478 = _T_2477 | _T_2463; // @[Mux.scala 27:72]
  wire  _T_2431 = _T_2409 == 4'h7; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2464 = _T_2431 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2479 = _T_2478 | _T_2464; // @[Mux.scala 27:72]
  wire  _T_2434 = _T_2409 == 4'h8; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2465 = _T_2434 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2480 = _T_2479 | _T_2465; // @[Mux.scala 27:72]
  wire  _T_2437 = _T_2409 == 4'h9; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2466 = _T_2437 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2481 = _T_2480 | _T_2466; // @[Mux.scala 27:72]
  wire  _T_2440 = _T_2409 == 4'ha; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2467 = _T_2440 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2482 = _T_2481 | _T_2467; // @[Mux.scala 27:72]
  wire  _T_2443 = _T_2409 == 4'hb; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2468 = _T_2443 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2483 = _T_2482 | _T_2468; // @[Mux.scala 27:72]
  wire  _T_2446 = _T_2409 == 4'hc; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2469 = _T_2446 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2484 = _T_2483 | _T_2469; // @[Mux.scala 27:72]
  wire  _T_2449 = _T_2409 == 4'hd; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2470 = _T_2449 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2485 = _T_2484 | _T_2470; // @[Mux.scala 27:72]
  wire  _T_2452 = _T_2409 == 4'he; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2471 = _T_2452 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2486 = _T_2485 | _T_2471; // @[Mux.scala 27:72]
  wire  _T_2455 = _T_2409 == 4'hf; // @[el2_ifu_mem_ctl.scala 475:66]
  wire [31:0] _T_2472 = _T_2455 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2487 = _T_2486 | _T_2472; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2407,_T_2487}; // @[Cat.scala 29:58]
  wire [6:0] _T_991 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 416:13]
  wire  _T_992 = ^_T_991; // @[el2_lib.scala 416:20]
  wire [6:0] _T_998 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_1005 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 416:30]
  wire [14:0] _T_1006 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_998}; // @[el2_lib.scala 416:30]
  wire [7:0] _T_1013 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 416:30]
  wire [30:0] _T_1022 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1013,_T_1006}; // @[el2_lib.scala 416:30]
  wire  _T_1023 = ^_T_1022; // @[el2_lib.scala 416:37]
  wire [6:0] _T_1029 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 416:47]
  wire [14:0] _T_1037 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1029}; // @[el2_lib.scala 416:47]
  wire [30:0] _T_1053 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1013,_T_1037}; // @[el2_lib.scala 416:47]
  wire  _T_1054 = ^_T_1053; // @[el2_lib.scala 416:54]
  wire [6:0] _T_1060 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 416:64]
  wire [14:0] _T_1068 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1060}; // @[el2_lib.scala 416:64]
  wire [30:0] _T_1084 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1005,_T_1068}; // @[el2_lib.scala 416:64]
  wire  _T_1085 = ^_T_1084; // @[el2_lib.scala 416:71]
  wire [7:0] _T_1092 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 416:81]
  wire [16:0] _T_1101 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1092}; // @[el2_lib.scala 416:81]
  wire [8:0] _T_1109 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 416:81]
  wire [17:0] _T_1118 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1109}; // @[el2_lib.scala 416:81]
  wire [34:0] _T_1119 = {_T_1118,_T_1101}; // @[el2_lib.scala 416:81]
  wire  _T_1120 = ^_T_1119; // @[el2_lib.scala 416:88]
  wire [7:0] _T_1127 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 416:98]
  wire [16:0] _T_1136 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1127}; // @[el2_lib.scala 416:98]
  wire [8:0] _T_1144 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 416:98]
  wire [17:0] _T_1153 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1144}; // @[el2_lib.scala 416:98]
  wire [34:0] _T_1154 = {_T_1153,_T_1136}; // @[el2_lib.scala 416:98]
  wire  _T_1155 = ^_T_1154; // @[el2_lib.scala 416:105]
  wire [7:0] _T_1162 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 416:115]
  wire [16:0] _T_1171 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_1162}; // @[el2_lib.scala 416:115]
  wire [8:0] _T_1179 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 416:115]
  wire [17:0] _T_1188 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1179}; // @[el2_lib.scala 416:115]
  wire [34:0] _T_1189 = {_T_1188,_T_1171}; // @[el2_lib.scala 416:115]
  wire  _T_1190 = ^_T_1189; // @[el2_lib.scala 416:122]
  wire [70:0] _T_1235 = {_T_570,_T_601,_T_632,_T_663,_T_698,_T_733,_T_768,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1234 = {_T_992,_T_1023,_T_1054,_T_1085,_T_1120,_T_1155,_T_1190,_T_2407,_T_2487}; // @[Cat.scala 29:58]
  wire [141:0] _T_1236 = {_T_570,_T_601,_T_632,_T_663,_T_698,_T_733,_T_768,ifu_bus_rdata_ff,_T_1234}; // @[Cat.scala 29:58]
  wire [141:0] _T_1239 = {_T_992,_T_1023,_T_1054,_T_1085,_T_1120,_T_1155,_T_1190,_T_2407,_T_2487,_T_1235}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1236 : _T_1239; // @[el2_ifu_mem_ctl.scala 359:28]
  wire  _T_1198 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 349:56]
  wire  _T_1199 = _T_1198 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 349:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 420:28]
  wire  _T_1403 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 422:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 624:35]
  wire  _T_1288 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 404:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 404:73]
  wire  _T_1329 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 411:118]
  wire  _T_1330 = ic_miss_buff_data_valid[0] & _T_1329; // @[el2_ifu_mem_ctl.scala 411:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1330; // @[el2_ifu_mem_ctl.scala 411:88]
  wire  _T_1426 = _T_1403 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1406 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 422:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 404:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 404:73]
  wire  _T_1333 = ic_miss_buff_data_valid[1] & _T_1329; // @[el2_ifu_mem_ctl.scala 411:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1333; // @[el2_ifu_mem_ctl.scala 411:88]
  wire  _T_1427 = _T_1406 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1434 = _T_1426 | _T_1427; // @[Mux.scala 27:72]
  wire  _T_1409 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 422:114]
  wire  _T_1290 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 404:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1290; // @[el2_ifu_mem_ctl.scala 404:73]
  wire  _T_1336 = ic_miss_buff_data_valid[2] & _T_1329; // @[el2_ifu_mem_ctl.scala 411:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1336; // @[el2_ifu_mem_ctl.scala 411:88]
  wire  _T_1428 = _T_1409 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1435 = _T_1434 | _T_1428; // @[Mux.scala 27:72]
  wire  _T_1412 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 422:114]
  wire  _T_1291 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 404:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1291; // @[el2_ifu_mem_ctl.scala 404:73]
  wire  _T_1339 = ic_miss_buff_data_valid[3] & _T_1329; // @[el2_ifu_mem_ctl.scala 411:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1339; // @[el2_ifu_mem_ctl.scala 411:88]
  wire  _T_1429 = _T_1412 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1436 = _T_1435 | _T_1429; // @[Mux.scala 27:72]
  wire  _T_1415 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 422:114]
  wire  _T_1292 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 404:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1292; // @[el2_ifu_mem_ctl.scala 404:73]
  wire  _T_1342 = ic_miss_buff_data_valid[4] & _T_1329; // @[el2_ifu_mem_ctl.scala 411:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1342; // @[el2_ifu_mem_ctl.scala 411:88]
  wire  _T_1430 = _T_1415 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1437 = _T_1436 | _T_1430; // @[Mux.scala 27:72]
  wire  _T_1418 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 422:114]
  wire  _T_1293 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 404:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1293; // @[el2_ifu_mem_ctl.scala 404:73]
  wire  _T_1345 = ic_miss_buff_data_valid[5] & _T_1329; // @[el2_ifu_mem_ctl.scala 411:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1345; // @[el2_ifu_mem_ctl.scala 411:88]
  wire  _T_1431 = _T_1418 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1438 = _T_1437 | _T_1431; // @[Mux.scala 27:72]
  wire  _T_1421 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 422:114]
  wire  _T_1294 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 404:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1294; // @[el2_ifu_mem_ctl.scala 404:73]
  wire  _T_1348 = ic_miss_buff_data_valid[6] & _T_1329; // @[el2_ifu_mem_ctl.scala 411:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1348; // @[el2_ifu_mem_ctl.scala 411:88]
  wire  _T_1432 = _T_1421 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1439 = _T_1438 | _T_1432; // @[Mux.scala 27:72]
  wire  _T_1424 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 422:114]
  wire  _T_1295 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 404:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1295; // @[el2_ifu_mem_ctl.scala 404:73]
  wire  _T_1351 = ic_miss_buff_data_valid[7] & _T_1329; // @[el2_ifu_mem_ctl.scala 411:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1351; // @[el2_ifu_mem_ctl.scala 411:88]
  wire  _T_1433 = _T_1424 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1439 | _T_1433; // @[Mux.scala 27:72]
  wire  _T_1442 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 423:58]
  wire  _T_1443 = bypass_valid_value_check & _T_1442; // @[el2_ifu_mem_ctl.scala 423:56]
  wire  _T_1445 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 423:77]
  wire  _T_1446 = _T_1443 & _T_1445; // @[el2_ifu_mem_ctl.scala 423:75]
  wire  _T_1451 = _T_1443 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 424:75]
  wire  _T_1452 = _T_1446 | _T_1451; // @[el2_ifu_mem_ctl.scala 423:95]
  wire  _T_1454 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 425:56]
  wire  _T_1457 = _T_1454 & _T_1445; // @[el2_ifu_mem_ctl.scala 425:74]
  wire  _T_1458 = _T_1452 | _T_1457; // @[el2_ifu_mem_ctl.scala 424:94]
  wire  _T_1462 = _T_1454 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 426:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 421:70]
  wire  _T_1463 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 426:132]
  wire  _T_1479 = _T_1463 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1465 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 426:132]
  wire  _T_1480 = _T_1465 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1487 = _T_1479 | _T_1480; // @[Mux.scala 27:72]
  wire  _T_1467 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 426:132]
  wire  _T_1481 = _T_1467 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1488 = _T_1487 | _T_1481; // @[Mux.scala 27:72]
  wire  _T_1469 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 426:132]
  wire  _T_1482 = _T_1469 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1489 = _T_1488 | _T_1482; // @[Mux.scala 27:72]
  wire  _T_1471 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 426:132]
  wire  _T_1483 = _T_1471 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1490 = _T_1489 | _T_1483; // @[Mux.scala 27:72]
  wire  _T_1473 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 426:132]
  wire  _T_1484 = _T_1473 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1491 = _T_1490 | _T_1484; // @[Mux.scala 27:72]
  wire  _T_1475 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 426:132]
  wire  _T_1485 = _T_1475 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1492 = _T_1491 | _T_1485; // @[Mux.scala 27:72]
  wire  _T_1477 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 426:132]
  wire  _T_1486 = _T_1477 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1493 = _T_1492 | _T_1486; // @[Mux.scala 27:72]
  wire  _T_1495 = _T_1462 & _T_1493; // @[el2_ifu_mem_ctl.scala 426:69]
  wire  _T_1496 = _T_1458 | _T_1495; // @[el2_ifu_mem_ctl.scala 425:94]
  wire [4:0] _GEN_437 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 427:95]
  wire  _T_1499 = _GEN_437 == 5'h1f; // @[el2_ifu_mem_ctl.scala 427:95]
  wire  _T_1500 = bypass_valid_value_check & _T_1499; // @[el2_ifu_mem_ctl.scala 427:56]
  wire  bypass_data_ready_in = _T_1496 | _T_1500; // @[el2_ifu_mem_ctl.scala 426:181]
  wire  _T_1501 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 431:53]
  wire  _T_1502 = _T_1501 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 431:73]
  wire  _T_1504 = _T_1502 & _T_319; // @[el2_ifu_mem_ctl.scala 431:96]
  wire  _T_1506 = _T_1504 & _T_58; // @[el2_ifu_mem_ctl.scala 431:118]
  wire  _T_1508 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 432:73]
  wire  _T_1510 = _T_1508 & _T_319; // @[el2_ifu_mem_ctl.scala 432:96]
  wire  _T_1512 = _T_1510 & _T_58; // @[el2_ifu_mem_ctl.scala 432:118]
  wire  _T_1513 = _T_1506 | _T_1512; // @[el2_ifu_mem_ctl.scala 431:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 434:58]
  wire  _T_1514 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 433:54]
  wire  _T_1515 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 433:76]
  wire  _T_1516 = _T_1514 & _T_1515; // @[el2_ifu_mem_ctl.scala 433:74]
  wire  _T_1518 = _T_1516 & _T_319; // @[el2_ifu_mem_ctl.scala 433:96]
  wire  ic_crit_wd_rdy_new_in = _T_1513 | _T_1518; // @[el2_ifu_mem_ctl.scala 432:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 634:43]
  wire  _T_1251 = ic_crit_wd_rdy | _T_2267; // @[el2_ifu_mem_ctl.scala 372:38]
  wire  _T_1253 = _T_1251 | _T_2283; // @[el2_ifu_mem_ctl.scala 372:64]
  wire  _T_1254 = ~_T_1253; // @[el2_ifu_mem_ctl.scala 372:21]
  wire  _T_1255 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 372:98]
  wire  sel_ic_data = _T_1254 & _T_1255; // @[el2_ifu_mem_ctl.scala 372:96]
  wire  _T_2490 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 477:44]
  wire  _T_1611 = ~ifu_fetch_addr_int_f[1]; // @[el2_ifu_mem_ctl.scala 444:30]
  wire  _T_1613 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 444:57]
  wire  _T_1614 = _T_1611 & _T_1613; // @[el2_ifu_mem_ctl.scala 444:55]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 417:60]
  wire [7:0] _T_1616 = ic_miss_buff_data_error >> byp_fetch_index[4:2]; // @[el2_ifu_mem_ctl.scala 444:107]
  wire  _T_1618 = _T_1614 & _T_1616[0]; // @[el2_ifu_mem_ctl.scala 444:82]
  wire  _T_1622 = _T_1611 & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 445:33]
  wire  _T_1626 = _T_1622 & _T_1616[0]; // @[el2_ifu_mem_ctl.scala 445:60]
  wire  _T_1627 = _T_1618 | _T_1626; // @[el2_ifu_mem_ctl.scala 444:151]
  wire  _T_1636 = _T_1627 | _T_1626; // @[el2_ifu_mem_ctl.scala 445:129]
  wire  _T_1640 = ifu_fetch_addr_int_f[1] & _T_1613; // @[el2_ifu_mem_ctl.scala 447:33]
  wire  _T_1644 = _T_1640 & _T_1616[0]; // @[el2_ifu_mem_ctl.scala 447:60]
  wire  _T_1645 = _T_1636 | _T_1644; // @[el2_ifu_mem_ctl.scala 446:129]
  wire  _T_1648 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 448:32]
  wire [7:0] _T_1653 = ic_miss_buff_data_error >> byp_fetch_index_inc; // @[el2_ifu_mem_ctl.scala 449:32]
  wire  _T_1655 = _T_1616[0] | _T_1653[0]; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_1656 = _T_1648 & _T_1655; // @[el2_ifu_mem_ctl.scala 448:58]
  wire  ifu_byp_data_err_new = _T_1645 | _T_1656; // @[el2_ifu_mem_ctl.scala 447:129]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 389:42]
  wire  _T_2491 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 477:91]
  wire  _T_2492 = ~_T_2491; // @[el2_ifu_mem_ctl.scala 477:60]
  wire  ic_rd_parity_final_err = _T_2490 & _T_2492; // @[el2_ifu_mem_ctl.scala 477:58]
  reg  ic_debug_ict_array_sel_ff; // @[el2_ifu_mem_ctl.scala 842:63]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9373 = _T_4670 & ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 769:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9375 = _T_4671 & ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9628 = _T_9373 | _T_9375; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9377 = _T_4672 & ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9629 = _T_9628 | _T_9377; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9379 = _T_4673 & ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9630 = _T_9629 | _T_9379; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9381 = _T_4674 & ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9631 = _T_9630 | _T_9381; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9383 = _T_4675 & ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9632 = _T_9631 | _T_9383; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9385 = _T_4676 & ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9633 = _T_9632 | _T_9385; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9387 = _T_4677 & ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9634 = _T_9633 | _T_9387; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9389 = _T_4678 & ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9635 = _T_9634 | _T_9389; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9391 = _T_4679 & ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9636 = _T_9635 | _T_9391; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9393 = _T_4680 & ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9637 = _T_9636 | _T_9393; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9395 = _T_4681 & ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9638 = _T_9637 | _T_9395; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9397 = _T_4682 & ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9639 = _T_9638 | _T_9397; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9399 = _T_4683 & ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9640 = _T_9639 | _T_9399; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9401 = _T_4684 & ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9641 = _T_9640 | _T_9401; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9403 = _T_4685 & ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9642 = _T_9641 | _T_9403; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9405 = _T_4686 & ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9643 = _T_9642 | _T_9405; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9407 = _T_4687 & ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9644 = _T_9643 | _T_9407; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9409 = _T_4688 & ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9645 = _T_9644 | _T_9409; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9411 = _T_4689 & ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9646 = _T_9645 | _T_9411; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9413 = _T_4690 & ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9647 = _T_9646 | _T_9413; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9415 = _T_4691 & ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9648 = _T_9647 | _T_9415; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9417 = _T_4692 & ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9649 = _T_9648 | _T_9417; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9419 = _T_4693 & ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9650 = _T_9649 | _T_9419; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9421 = _T_4694 & ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9651 = _T_9650 | _T_9421; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9423 = _T_4695 & ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9652 = _T_9651 | _T_9423; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9425 = _T_4696 & ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9653 = _T_9652 | _T_9425; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9427 = _T_4697 & ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9654 = _T_9653 | _T_9427; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9429 = _T_4698 & ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9655 = _T_9654 | _T_9429; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9431 = _T_4699 & ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9656 = _T_9655 | _T_9431; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9433 = _T_4700 & ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9657 = _T_9656 | _T_9433; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9435 = _T_4701 & ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9658 = _T_9657 | _T_9435; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9437 = _T_4702 & ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9659 = _T_9658 | _T_9437; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9439 = _T_4703 & ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9660 = _T_9659 | _T_9439; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9441 = _T_4704 & ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9661 = _T_9660 | _T_9441; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9443 = _T_4705 & ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9662 = _T_9661 | _T_9443; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9445 = _T_4706 & ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9663 = _T_9662 | _T_9445; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9447 = _T_4707 & ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9664 = _T_9663 | _T_9447; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9449 = _T_4708 & ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9665 = _T_9664 | _T_9449; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9451 = _T_4709 & ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9666 = _T_9665 | _T_9451; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9453 = _T_4710 & ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9667 = _T_9666 | _T_9453; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9455 = _T_4711 & ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9668 = _T_9667 | _T_9455; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9457 = _T_4712 & ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9669 = _T_9668 | _T_9457; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9459 = _T_4713 & ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9670 = _T_9669 | _T_9459; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9461 = _T_4714 & ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9671 = _T_9670 | _T_9461; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9463 = _T_4715 & ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9672 = _T_9671 | _T_9463; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9465 = _T_4716 & ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9673 = _T_9672 | _T_9465; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9467 = _T_4717 & ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9674 = _T_9673 | _T_9467; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9469 = _T_4718 & ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9675 = _T_9674 | _T_9469; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9471 = _T_4719 & ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9676 = _T_9675 | _T_9471; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9473 = _T_4720 & ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9677 = _T_9676 | _T_9473; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9475 = _T_4721 & ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9678 = _T_9677 | _T_9475; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9477 = _T_4722 & ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9679 = _T_9678 | _T_9477; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9479 = _T_4723 & ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9680 = _T_9679 | _T_9479; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9481 = _T_4724 & ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9681 = _T_9680 | _T_9481; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9483 = _T_4725 & ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9682 = _T_9681 | _T_9483; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9485 = _T_4726 & ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9683 = _T_9682 | _T_9485; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9487 = _T_4727 & ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9684 = _T_9683 | _T_9487; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9489 = _T_4728 & ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9685 = _T_9684 | _T_9489; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9491 = _T_4729 & ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9686 = _T_9685 | _T_9491; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9493 = _T_4730 & ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9687 = _T_9686 | _T_9493; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9495 = _T_4731 & ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9688 = _T_9687 | _T_9495; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9497 = _T_4732 & ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9689 = _T_9688 | _T_9497; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9499 = _T_4733 & ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9690 = _T_9689 | _T_9499; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9501 = _T_4734 & ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9691 = _T_9690 | _T_9501; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9503 = _T_4735 & ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9692 = _T_9691 | _T_9503; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9505 = _T_4736 & ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9693 = _T_9692 | _T_9505; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9507 = _T_4737 & ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9694 = _T_9693 | _T_9507; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9509 = _T_4738 & ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9695 = _T_9694 | _T_9509; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9511 = _T_4739 & ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9696 = _T_9695 | _T_9511; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9513 = _T_4740 & ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9697 = _T_9696 | _T_9513; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9515 = _T_4741 & ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9698 = _T_9697 | _T_9515; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9517 = _T_4742 & ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9699 = _T_9698 | _T_9517; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9519 = _T_4743 & ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9700 = _T_9699 | _T_9519; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9521 = _T_4744 & ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9701 = _T_9700 | _T_9521; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9523 = _T_4745 & ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9702 = _T_9701 | _T_9523; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9525 = _T_4746 & ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9703 = _T_9702 | _T_9525; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9527 = _T_4747 & ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9704 = _T_9703 | _T_9527; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9529 = _T_4748 & ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9705 = _T_9704 | _T_9529; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9531 = _T_4749 & ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9706 = _T_9705 | _T_9531; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9533 = _T_4750 & ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9707 = _T_9706 | _T_9533; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9535 = _T_4751 & ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9708 = _T_9707 | _T_9535; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9537 = _T_4752 & ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9709 = _T_9708 | _T_9537; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9539 = _T_4753 & ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9710 = _T_9709 | _T_9539; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9541 = _T_4754 & ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9711 = _T_9710 | _T_9541; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9543 = _T_4755 & ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9712 = _T_9711 | _T_9543; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9545 = _T_4756 & ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9713 = _T_9712 | _T_9545; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9547 = _T_4757 & ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9714 = _T_9713 | _T_9547; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9549 = _T_4758 & ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9715 = _T_9714 | _T_9549; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9551 = _T_4759 & ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9716 = _T_9715 | _T_9551; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9553 = _T_4760 & ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9717 = _T_9716 | _T_9553; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9555 = _T_4761 & ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9718 = _T_9717 | _T_9555; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9557 = _T_4762 & ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9719 = _T_9718 | _T_9557; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9559 = _T_4763 & ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9720 = _T_9719 | _T_9559; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9561 = _T_4764 & ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9721 = _T_9720 | _T_9561; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9563 = _T_4765 & ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9722 = _T_9721 | _T_9563; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9565 = _T_4766 & ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9723 = _T_9722 | _T_9565; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9567 = _T_4767 & ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9724 = _T_9723 | _T_9567; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9569 = _T_4768 & ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9725 = _T_9724 | _T_9569; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9571 = _T_4769 & ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9726 = _T_9725 | _T_9571; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9573 = _T_4770 & ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9727 = _T_9726 | _T_9573; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9575 = _T_4771 & ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9728 = _T_9727 | _T_9575; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9577 = _T_4772 & ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9729 = _T_9728 | _T_9577; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9579 = _T_4773 & ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9730 = _T_9729 | _T_9579; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9581 = _T_4774 & ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9731 = _T_9730 | _T_9581; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9583 = _T_4775 & ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9732 = _T_9731 | _T_9583; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9585 = _T_4776 & ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9733 = _T_9732 | _T_9585; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9587 = _T_4777 & ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9734 = _T_9733 | _T_9587; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9589 = _T_4778 & ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9735 = _T_9734 | _T_9589; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9591 = _T_4779 & ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9736 = _T_9735 | _T_9591; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9593 = _T_4780 & ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9737 = _T_9736 | _T_9593; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9595 = _T_4781 & ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9738 = _T_9737 | _T_9595; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9597 = _T_4782 & ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9739 = _T_9738 | _T_9597; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9599 = _T_4783 & ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9740 = _T_9739 | _T_9599; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9601 = _T_4784 & ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9741 = _T_9740 | _T_9601; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9603 = _T_4785 & ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9742 = _T_9741 | _T_9603; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9605 = _T_4786 & ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9743 = _T_9742 | _T_9605; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9607 = _T_4787 & ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9744 = _T_9743 | _T_9607; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9609 = _T_4788 & ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9745 = _T_9744 | _T_9609; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9611 = _T_4789 & ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9746 = _T_9745 | _T_9611; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9613 = _T_4790 & ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9747 = _T_9746 | _T_9613; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9615 = _T_4791 & ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9748 = _T_9747 | _T_9615; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9617 = _T_4792 & ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9749 = _T_9748 | _T_9617; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9619 = _T_4793 & ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9750 = _T_9749 | _T_9619; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9621 = _T_4794 & ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9751 = _T_9750 | _T_9621; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9623 = _T_4795 & ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9752 = _T_9751 | _T_9623; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9625 = _T_4796 & ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9753 = _T_9752 | _T_9625; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9627 = _T_4797 & ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9754 = _T_9753 | _T_9627; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_8990 = _T_4670 & ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 769:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_8992 = _T_4671 & ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9245 = _T_8990 | _T_8992; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_8994 = _T_4672 & ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9246 = _T_9245 | _T_8994; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_8996 = _T_4673 & ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9247 = _T_9246 | _T_8996; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_8998 = _T_4674 & ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9248 = _T_9247 | _T_8998; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9000 = _T_4675 & ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9249 = _T_9248 | _T_9000; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9002 = _T_4676 & ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9250 = _T_9249 | _T_9002; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9004 = _T_4677 & ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9251 = _T_9250 | _T_9004; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9006 = _T_4678 & ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9252 = _T_9251 | _T_9006; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9008 = _T_4679 & ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9253 = _T_9252 | _T_9008; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9010 = _T_4680 & ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9254 = _T_9253 | _T_9010; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9012 = _T_4681 & ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9255 = _T_9254 | _T_9012; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9014 = _T_4682 & ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9256 = _T_9255 | _T_9014; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9016 = _T_4683 & ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9257 = _T_9256 | _T_9016; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9018 = _T_4684 & ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9258 = _T_9257 | _T_9018; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9020 = _T_4685 & ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9259 = _T_9258 | _T_9020; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9022 = _T_4686 & ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9260 = _T_9259 | _T_9022; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9024 = _T_4687 & ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9261 = _T_9260 | _T_9024; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9026 = _T_4688 & ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9262 = _T_9261 | _T_9026; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9028 = _T_4689 & ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9263 = _T_9262 | _T_9028; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9030 = _T_4690 & ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9264 = _T_9263 | _T_9030; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9032 = _T_4691 & ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9265 = _T_9264 | _T_9032; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9034 = _T_4692 & ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9266 = _T_9265 | _T_9034; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9036 = _T_4693 & ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9267 = _T_9266 | _T_9036; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9038 = _T_4694 & ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9268 = _T_9267 | _T_9038; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9040 = _T_4695 & ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9269 = _T_9268 | _T_9040; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9042 = _T_4696 & ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9270 = _T_9269 | _T_9042; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9044 = _T_4697 & ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9271 = _T_9270 | _T_9044; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9046 = _T_4698 & ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9272 = _T_9271 | _T_9046; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9048 = _T_4699 & ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9273 = _T_9272 | _T_9048; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9050 = _T_4700 & ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9274 = _T_9273 | _T_9050; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9052 = _T_4701 & ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9275 = _T_9274 | _T_9052; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9054 = _T_4702 & ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9276 = _T_9275 | _T_9054; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9056 = _T_4703 & ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9277 = _T_9276 | _T_9056; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9058 = _T_4704 & ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9278 = _T_9277 | _T_9058; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9060 = _T_4705 & ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9279 = _T_9278 | _T_9060; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9062 = _T_4706 & ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9280 = _T_9279 | _T_9062; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9064 = _T_4707 & ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9281 = _T_9280 | _T_9064; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9066 = _T_4708 & ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9282 = _T_9281 | _T_9066; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9068 = _T_4709 & ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9283 = _T_9282 | _T_9068; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9070 = _T_4710 & ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9284 = _T_9283 | _T_9070; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9072 = _T_4711 & ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9285 = _T_9284 | _T_9072; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9074 = _T_4712 & ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9286 = _T_9285 | _T_9074; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9076 = _T_4713 & ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9287 = _T_9286 | _T_9076; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9078 = _T_4714 & ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9288 = _T_9287 | _T_9078; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9080 = _T_4715 & ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9289 = _T_9288 | _T_9080; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9082 = _T_4716 & ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9290 = _T_9289 | _T_9082; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9084 = _T_4717 & ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9291 = _T_9290 | _T_9084; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9086 = _T_4718 & ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9292 = _T_9291 | _T_9086; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9088 = _T_4719 & ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9293 = _T_9292 | _T_9088; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9090 = _T_4720 & ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9294 = _T_9293 | _T_9090; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9092 = _T_4721 & ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9295 = _T_9294 | _T_9092; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9094 = _T_4722 & ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9296 = _T_9295 | _T_9094; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9096 = _T_4723 & ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9297 = _T_9296 | _T_9096; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9098 = _T_4724 & ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9298 = _T_9297 | _T_9098; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9100 = _T_4725 & ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9299 = _T_9298 | _T_9100; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9102 = _T_4726 & ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9300 = _T_9299 | _T_9102; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9104 = _T_4727 & ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9301 = _T_9300 | _T_9104; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9106 = _T_4728 & ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9302 = _T_9301 | _T_9106; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9108 = _T_4729 & ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9303 = _T_9302 | _T_9108; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9110 = _T_4730 & ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9304 = _T_9303 | _T_9110; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9112 = _T_4731 & ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9305 = _T_9304 | _T_9112; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9114 = _T_4732 & ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9306 = _T_9305 | _T_9114; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9116 = _T_4733 & ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9307 = _T_9306 | _T_9116; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9118 = _T_4734 & ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9308 = _T_9307 | _T_9118; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9120 = _T_4735 & ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9309 = _T_9308 | _T_9120; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9122 = _T_4736 & ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9310 = _T_9309 | _T_9122; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9124 = _T_4737 & ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9311 = _T_9310 | _T_9124; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9126 = _T_4738 & ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9312 = _T_9311 | _T_9126; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9128 = _T_4739 & ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9313 = _T_9312 | _T_9128; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9130 = _T_4740 & ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9314 = _T_9313 | _T_9130; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9132 = _T_4741 & ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9315 = _T_9314 | _T_9132; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9134 = _T_4742 & ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9316 = _T_9315 | _T_9134; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9136 = _T_4743 & ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9317 = _T_9316 | _T_9136; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9138 = _T_4744 & ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9318 = _T_9317 | _T_9138; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9140 = _T_4745 & ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9319 = _T_9318 | _T_9140; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9142 = _T_4746 & ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9320 = _T_9319 | _T_9142; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9144 = _T_4747 & ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9321 = _T_9320 | _T_9144; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9146 = _T_4748 & ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9322 = _T_9321 | _T_9146; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9148 = _T_4749 & ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9323 = _T_9322 | _T_9148; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9150 = _T_4750 & ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9324 = _T_9323 | _T_9150; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9152 = _T_4751 & ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9325 = _T_9324 | _T_9152; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9154 = _T_4752 & ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9326 = _T_9325 | _T_9154; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9156 = _T_4753 & ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9327 = _T_9326 | _T_9156; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9158 = _T_4754 & ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9328 = _T_9327 | _T_9158; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9160 = _T_4755 & ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9329 = _T_9328 | _T_9160; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9162 = _T_4756 & ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9330 = _T_9329 | _T_9162; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9164 = _T_4757 & ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9331 = _T_9330 | _T_9164; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9166 = _T_4758 & ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9332 = _T_9331 | _T_9166; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9168 = _T_4759 & ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9333 = _T_9332 | _T_9168; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9170 = _T_4760 & ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9334 = _T_9333 | _T_9170; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9172 = _T_4761 & ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9335 = _T_9334 | _T_9172; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9174 = _T_4762 & ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9336 = _T_9335 | _T_9174; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9176 = _T_4763 & ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9337 = _T_9336 | _T_9176; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9178 = _T_4764 & ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9338 = _T_9337 | _T_9178; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9180 = _T_4765 & ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9339 = _T_9338 | _T_9180; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9182 = _T_4766 & ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9340 = _T_9339 | _T_9182; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9184 = _T_4767 & ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9341 = _T_9340 | _T_9184; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9186 = _T_4768 & ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9342 = _T_9341 | _T_9186; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9188 = _T_4769 & ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9343 = _T_9342 | _T_9188; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9190 = _T_4770 & ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9344 = _T_9343 | _T_9190; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9192 = _T_4771 & ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9345 = _T_9344 | _T_9192; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9194 = _T_4772 & ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9346 = _T_9345 | _T_9194; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9196 = _T_4773 & ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9347 = _T_9346 | _T_9196; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9198 = _T_4774 & ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9348 = _T_9347 | _T_9198; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9200 = _T_4775 & ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9349 = _T_9348 | _T_9200; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9202 = _T_4776 & ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9350 = _T_9349 | _T_9202; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9204 = _T_4777 & ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9351 = _T_9350 | _T_9204; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9206 = _T_4778 & ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9352 = _T_9351 | _T_9206; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9208 = _T_4779 & ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9353 = _T_9352 | _T_9208; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9210 = _T_4780 & ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9354 = _T_9353 | _T_9210; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9212 = _T_4781 & ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9355 = _T_9354 | _T_9212; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9214 = _T_4782 & ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9356 = _T_9355 | _T_9214; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9216 = _T_4783 & ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9357 = _T_9356 | _T_9216; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9218 = _T_4784 & ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9358 = _T_9357 | _T_9218; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9220 = _T_4785 & ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9359 = _T_9358 | _T_9220; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9222 = _T_4786 & ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9360 = _T_9359 | _T_9222; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9224 = _T_4787 & ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9361 = _T_9360 | _T_9224; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9226 = _T_4788 & ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9362 = _T_9361 | _T_9226; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9228 = _T_4789 & ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9363 = _T_9362 | _T_9228; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9230 = _T_4790 & ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9364 = _T_9363 | _T_9230; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9232 = _T_4791 & ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9365 = _T_9364 | _T_9232; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9234 = _T_4792 & ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9366 = _T_9365 | _T_9234; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9236 = _T_4793 & ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9367 = _T_9366 | _T_9236; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9238 = _T_4794 & ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9368 = _T_9367 | _T_9238; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9240 = _T_4795 & ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9369 = _T_9368 | _T_9240; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9242 = _T_4796 & ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9370 = _T_9369 | _T_9242; // @[el2_ifu_mem_ctl.scala 769:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9244 = _T_4797 & ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 769:10]
  wire  _T_9371 = _T_9370 | _T_9244; // @[el2_ifu_mem_ctl.scala 769:91]
  wire [1:0] ic_tag_valid_unq = {_T_9754,_T_9371}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[el2_ifu_mem_ctl.scala 841:53]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 843:54]
  wire [1:0] _T_9794 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_9795 = ic_debug_way_ff & _T_9794; // @[el2_ifu_mem_ctl.scala 824:67]
  wire [1:0] _T_9796 = ic_tag_valid_unq & _T_9795; // @[el2_ifu_mem_ctl.scala 824:48]
  wire  ic_debug_tag_val_rd_out = |_T_9796; // @[el2_ifu_mem_ctl.scala 824:115]
  wire [70:0] _T_1210 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],6'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1211; // @[el2_ifu_mem_ctl.scala 355:63]
  wire  _T_1249 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 371:98]
  wire  sel_byp_data = _T_1253 & _T_1249; // @[el2_ifu_mem_ctl.scala 371:96]
  wire  _T_1256 = sel_byp_data | fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 376:46]
  wire  final_data_sel1_0 = _T_1256 | sel_ic_data; // @[el2_ifu_mem_ctl.scala 376:62]
  wire [63:0] _T_1262 = final_data_sel1_0 ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] ic_final_data = _T_1262 & io_ic_rd_data; // @[el2_ifu_mem_ctl.scala 380:92]
  wire [63:0] _T_1264 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1265 = _T_1264 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 384:69]
  wire [63:0] _T_1267 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1661 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1709 = _T_1661 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1664 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1710 = _T_1664 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1725 = _T_1709 | _T_1710; // @[Mux.scala 27:72]
  wire  _T_1667 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1711 = _T_1667 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1726 = _T_1725 | _T_1711; // @[Mux.scala 27:72]
  wire  _T_1670 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1712 = _T_1670 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1727 = _T_1726 | _T_1712; // @[Mux.scala 27:72]
  wire  _T_1673 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1713 = _T_1673 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1728 = _T_1727 | _T_1713; // @[Mux.scala 27:72]
  wire  _T_1676 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1714 = _T_1676 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1729 = _T_1728 | _T_1714; // @[Mux.scala 27:72]
  wire  _T_1679 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1715 = _T_1679 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1730 = _T_1729 | _T_1715; // @[Mux.scala 27:72]
  wire  _T_1682 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1716 = _T_1682 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1731 = _T_1730 | _T_1716; // @[Mux.scala 27:72]
  wire  _T_1685 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1717 = _T_1685 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1732 = _T_1731 | _T_1717; // @[Mux.scala 27:72]
  wire  _T_1688 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1718 = _T_1688 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1733 = _T_1732 | _T_1718; // @[Mux.scala 27:72]
  wire  _T_1691 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1719 = _T_1691 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1734 = _T_1733 | _T_1719; // @[Mux.scala 27:72]
  wire  _T_1694 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1720 = _T_1694 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1735 = _T_1734 | _T_1720; // @[Mux.scala 27:72]
  wire  _T_1697 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1721 = _T_1697 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1736 = _T_1735 | _T_1721; // @[Mux.scala 27:72]
  wire  _T_1700 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1722 = _T_1700 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1737 = _T_1736 | _T_1722; // @[Mux.scala 27:72]
  wire  _T_1703 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1723 = _T_1703 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1738 = _T_1737 | _T_1723; // @[Mux.scala 27:72]
  wire  _T_1706 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 451:73]
  wire [15:0] _T_1724 = _T_1706 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1739 = _T_1738 | _T_1724; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1741 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1789 = _T_1741 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1744 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1790 = _T_1744 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1805 = _T_1789 | _T_1790; // @[Mux.scala 27:72]
  wire  _T_1747 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1791 = _T_1747 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1806 = _T_1805 | _T_1791; // @[Mux.scala 27:72]
  wire  _T_1750 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1792 = _T_1750 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1807 = _T_1806 | _T_1792; // @[Mux.scala 27:72]
  wire  _T_1753 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1793 = _T_1753 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1808 = _T_1807 | _T_1793; // @[Mux.scala 27:72]
  wire  _T_1756 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1794 = _T_1756 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1809 = _T_1808 | _T_1794; // @[Mux.scala 27:72]
  wire  _T_1759 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1795 = _T_1759 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1810 = _T_1809 | _T_1795; // @[Mux.scala 27:72]
  wire  _T_1762 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1796 = _T_1762 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1811 = _T_1810 | _T_1796; // @[Mux.scala 27:72]
  wire  _T_1765 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1797 = _T_1765 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1812 = _T_1811 | _T_1797; // @[Mux.scala 27:72]
  wire  _T_1768 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1798 = _T_1768 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1813 = _T_1812 | _T_1798; // @[Mux.scala 27:72]
  wire  _T_1771 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1799 = _T_1771 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1814 = _T_1813 | _T_1799; // @[Mux.scala 27:72]
  wire  _T_1774 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1800 = _T_1774 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1815 = _T_1814 | _T_1800; // @[Mux.scala 27:72]
  wire  _T_1777 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1801 = _T_1777 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1816 = _T_1815 | _T_1801; // @[Mux.scala 27:72]
  wire  _T_1780 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1802 = _T_1780 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1817 = _T_1816 | _T_1802; // @[Mux.scala 27:72]
  wire  _T_1783 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1803 = _T_1783 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1818 = _T_1817 | _T_1803; // @[Mux.scala 27:72]
  wire  _T_1786 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 451:179]
  wire [31:0] _T_1804 = _T_1786 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1819 = _T_1818 | _T_1804; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1821 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1869 = _T_1821 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1824 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1870 = _T_1824 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1885 = _T_1869 | _T_1870; // @[Mux.scala 27:72]
  wire  _T_1827 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1871 = _T_1827 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1886 = _T_1885 | _T_1871; // @[Mux.scala 27:72]
  wire  _T_1830 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1872 = _T_1830 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1887 = _T_1886 | _T_1872; // @[Mux.scala 27:72]
  wire  _T_1833 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1873 = _T_1833 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1888 = _T_1887 | _T_1873; // @[Mux.scala 27:72]
  wire  _T_1836 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1874 = _T_1836 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1889 = _T_1888 | _T_1874; // @[Mux.scala 27:72]
  wire  _T_1839 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1875 = _T_1839 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1890 = _T_1889 | _T_1875; // @[Mux.scala 27:72]
  wire  _T_1842 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1876 = _T_1842 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1891 = _T_1890 | _T_1876; // @[Mux.scala 27:72]
  wire  _T_1845 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1877 = _T_1845 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1892 = _T_1891 | _T_1877; // @[Mux.scala 27:72]
  wire  _T_1848 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1878 = _T_1848 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1893 = _T_1892 | _T_1878; // @[Mux.scala 27:72]
  wire  _T_1851 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1879 = _T_1851 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1894 = _T_1893 | _T_1879; // @[Mux.scala 27:72]
  wire  _T_1854 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1880 = _T_1854 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1895 = _T_1894 | _T_1880; // @[Mux.scala 27:72]
  wire  _T_1857 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1881 = _T_1857 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1896 = _T_1895 | _T_1881; // @[Mux.scala 27:72]
  wire  _T_1860 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1882 = _T_1860 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1897 = _T_1896 | _T_1882; // @[Mux.scala 27:72]
  wire  _T_1863 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1883 = _T_1863 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1898 = _T_1897 | _T_1883; // @[Mux.scala 27:72]
  wire  _T_1866 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 451:285]
  wire [31:0] _T_1884 = _T_1866 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1899 = _T_1898 | _T_1884; // @[Mux.scala 27:72]
  wire [79:0] _T_1902 = {_T_1739,_T_1819,_T_1899}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1903 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1951 = _T_1903 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1906 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1952 = _T_1906 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1967 = _T_1951 | _T_1952; // @[Mux.scala 27:72]
  wire  _T_1909 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1953 = _T_1909 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1968 = _T_1967 | _T_1953; // @[Mux.scala 27:72]
  wire  _T_1912 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1954 = _T_1912 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1969 = _T_1968 | _T_1954; // @[Mux.scala 27:72]
  wire  _T_1915 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1955 = _T_1915 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1970 = _T_1969 | _T_1955; // @[Mux.scala 27:72]
  wire  _T_1918 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1956 = _T_1918 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1971 = _T_1970 | _T_1956; // @[Mux.scala 27:72]
  wire  _T_1921 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1957 = _T_1921 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1972 = _T_1971 | _T_1957; // @[Mux.scala 27:72]
  wire  _T_1924 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1958 = _T_1924 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1973 = _T_1972 | _T_1958; // @[Mux.scala 27:72]
  wire  _T_1927 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1959 = _T_1927 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1974 = _T_1973 | _T_1959; // @[Mux.scala 27:72]
  wire  _T_1930 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1960 = _T_1930 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1975 = _T_1974 | _T_1960; // @[Mux.scala 27:72]
  wire  _T_1933 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1961 = _T_1933 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1976 = _T_1975 | _T_1961; // @[Mux.scala 27:72]
  wire  _T_1936 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1962 = _T_1936 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1977 = _T_1976 | _T_1962; // @[Mux.scala 27:72]
  wire  _T_1939 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1963 = _T_1939 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1978 = _T_1977 | _T_1963; // @[Mux.scala 27:72]
  wire  _T_1942 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1964 = _T_1942 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1979 = _T_1978 | _T_1964; // @[Mux.scala 27:72]
  wire  _T_1945 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1965 = _T_1945 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1980 = _T_1979 | _T_1965; // @[Mux.scala 27:72]
  wire  _T_1948 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_1966 = _T_1948 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1981 = _T_1980 | _T_1966; // @[Mux.scala 27:72]
  wire [31:0] _T_2031 = _T_1661 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2032 = _T_1664 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2047 = _T_2031 | _T_2032; // @[Mux.scala 27:72]
  wire [31:0] _T_2033 = _T_1667 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2048 = _T_2047 | _T_2033; // @[Mux.scala 27:72]
  wire [31:0] _T_2034 = _T_1670 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2049 = _T_2048 | _T_2034; // @[Mux.scala 27:72]
  wire [31:0] _T_2035 = _T_1673 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2050 = _T_2049 | _T_2035; // @[Mux.scala 27:72]
  wire [31:0] _T_2036 = _T_1676 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2051 = _T_2050 | _T_2036; // @[Mux.scala 27:72]
  wire [31:0] _T_2037 = _T_1679 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2052 = _T_2051 | _T_2037; // @[Mux.scala 27:72]
  wire [31:0] _T_2038 = _T_1682 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2053 = _T_2052 | _T_2038; // @[Mux.scala 27:72]
  wire [31:0] _T_2039 = _T_1685 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2054 = _T_2053 | _T_2039; // @[Mux.scala 27:72]
  wire [31:0] _T_2040 = _T_1688 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2055 = _T_2054 | _T_2040; // @[Mux.scala 27:72]
  wire [31:0] _T_2041 = _T_1691 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2056 = _T_2055 | _T_2041; // @[Mux.scala 27:72]
  wire [31:0] _T_2042 = _T_1694 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2057 = _T_2056 | _T_2042; // @[Mux.scala 27:72]
  wire [31:0] _T_2043 = _T_1697 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2058 = _T_2057 | _T_2043; // @[Mux.scala 27:72]
  wire [31:0] _T_2044 = _T_1700 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2059 = _T_2058 | _T_2044; // @[Mux.scala 27:72]
  wire [31:0] _T_2045 = _T_1703 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2060 = _T_2059 | _T_2045; // @[Mux.scala 27:72]
  wire [31:0] _T_2046 = _T_1706 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2061 = _T_2060 | _T_2046; // @[Mux.scala 27:72]
  wire [79:0] _T_2144 = {_T_1981,_T_2061,_T_1819}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1611 ? _T_1902 : _T_2144; // @[el2_ifu_mem_ctl.scala 450:37]
  wire [79:0] _T_2149 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_1613 ? ic_byp_data_only_pre_new : _T_2149; // @[el2_ifu_mem_ctl.scala 454:30]
  wire [79:0] _GEN_438 = {{16'd0}, _T_1267}; // @[el2_ifu_mem_ctl.scala 384:114]
  wire [79:0] _T_1268 = _GEN_438 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 384:114]
  wire [79:0] _GEN_439 = {{16'd0}, _T_1265}; // @[el2_ifu_mem_ctl.scala 384:88]
  wire [79:0] ic_premux_data_temp = _GEN_439 | _T_1268; // @[el2_ifu_mem_ctl.scala 384:88]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_319; // @[el2_ifu_mem_ctl.scala 391:38]
  reg  ifc_region_acc_fault_memory_f; // @[el2_ifu_mem_ctl.scala 856:66]
  wire [1:0] _T_1276 = ifc_region_acc_fault_memory_f ? 2'h3 : 2'h0; // @[el2_ifu_mem_ctl.scala 396:10]
  wire [1:0] _T_1277 = ifc_region_acc_fault_f ? 2'h2 : _T_1276; // @[el2_ifu_mem_ctl.scala 395:8]
  wire  _T_1279 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[el2_ifu_mem_ctl.scala 397:45]
  wire  _T_1281 = byp_fetch_index == 5'h1f; // @[el2_ifu_mem_ctl.scala 397:80]
  wire  _T_1282 = ~_T_1281; // @[el2_ifu_mem_ctl.scala 397:71]
  wire  _T_1283 = _T_1279 & _T_1282; // @[el2_ifu_mem_ctl.scala 397:69]
  wire  _T_1284 = err_stop_state != 2'h2; // @[el2_ifu_mem_ctl.scala 397:131]
  wire  _T_1285 = _T_1283 & _T_1284; // @[el2_ifu_mem_ctl.scala 397:114]
  wire [6:0] _T_1357 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1}; // @[Cat.scala 29:58]
  wire  _T_1363 = ic_miss_buff_data_error[0] & _T_1329; // @[el2_ifu_mem_ctl.scala 416:32]
  wire  _T_2689 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 630:47]
  wire  _T_2690 = _T_2689 & _T_13; // @[el2_ifu_mem_ctl.scala 630:50]
  wire  bus_ifu_wr_data_error = _T_2690 & miss_pending; // @[el2_ifu_mem_ctl.scala 630:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1363; // @[el2_ifu_mem_ctl.scala 415:72]
  wire  _T_1367 = ic_miss_buff_data_error[1] & _T_1329; // @[el2_ifu_mem_ctl.scala 416:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1367; // @[el2_ifu_mem_ctl.scala 415:72]
  wire  _T_1371 = ic_miss_buff_data_error[2] & _T_1329; // @[el2_ifu_mem_ctl.scala 416:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1371; // @[el2_ifu_mem_ctl.scala 415:72]
  wire  _T_1375 = ic_miss_buff_data_error[3] & _T_1329; // @[el2_ifu_mem_ctl.scala 416:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1375; // @[el2_ifu_mem_ctl.scala 415:72]
  wire  _T_1379 = ic_miss_buff_data_error[4] & _T_1329; // @[el2_ifu_mem_ctl.scala 416:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1379; // @[el2_ifu_mem_ctl.scala 415:72]
  wire  _T_1383 = ic_miss_buff_data_error[5] & _T_1329; // @[el2_ifu_mem_ctl.scala 416:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1383; // @[el2_ifu_mem_ctl.scala 415:72]
  wire  _T_1387 = ic_miss_buff_data_error[6] & _T_1329; // @[el2_ifu_mem_ctl.scala 416:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1387; // @[el2_ifu_mem_ctl.scala 415:72]
  wire  _T_1391 = ic_miss_buff_data_error[7] & _T_1329; // @[el2_ifu_mem_ctl.scala 416:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1391; // @[el2_ifu_mem_ctl.scala 415:72]
  wire [6:0] _T_1397 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1}; // @[Cat.scala 29:58]
  reg [6:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2499 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2507 = _T_6 & _T_319; // @[el2_ifu_mem_ctl.scala 497:65]
  wire  _T_2508 = _T_2507 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 497:88]
  wire  _T_2510 = _T_2508 & _T_2622; // @[el2_ifu_mem_ctl.scala 497:112]
  wire  _T_2511 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2512 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 502:50]
  wire  _T_2514 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2521 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2523 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_21 = _T_2521 | _T_2523; // @[Conditional.scala 39:67]
  wire  _GEN_23 = _T_2514 ? _T_2512 : _GEN_21; // @[Conditional.scala 39:67]
  wire  _GEN_25 = _T_2511 ? _T_2512 : _GEN_23; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2499 ? _T_2510 : _GEN_25; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2499 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2513 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 503:56]
  wire  _GEN_26 = _T_2511 & _T_2513; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2499 ? 1'h0 : _GEN_26; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 488:58]
  wire  _T_2496 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 487:49]
  wire  _T_2501 = io_ic_error_start & _T_319; // @[el2_ifu_mem_ctl.scala 496:87]
  wire  _T_2515 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 506:30]
  wire  _T_2516 = _T_2515 & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 506:55]
  wire  _T_2517 = _T_2516 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 506:85]
  wire  _T_2526 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 527:66]
  wire  _T_2527 = io_dec_tlu_flush_err_wb & _T_2526; // @[el2_ifu_mem_ctl.scala 527:52]
  wire  _T_2529 = _T_2527 & _T_2622; // @[el2_ifu_mem_ctl.scala 527:81]
  wire  _T_2531 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 530:59]
  wire  _T_2532 = _T_2531 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 530:86]
  wire  _T_2546 = _T_2531 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 533:81]
  wire  _T_2547 = _T_2546 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 533:103]
  wire  _T_2548 = _T_2547 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 533:126]
  wire  _T_2568 = _T_2546 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 540:103]
  wire  _T_2576 = io_dec_tlu_flush_lower_wb & _T_2515; // @[el2_ifu_mem_ctl.scala 545:60]
  wire  _T_2577 = _T_2576 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 545:88]
  wire  _T_2578 = _T_2577 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 545:115]
  wire  _GEN_33 = _T_2574 & _T_2532; // @[Conditional.scala 39:67]
  wire  _GEN_36 = _T_2557 ? _T_2568 : _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_38 = _T_2557 | _T_2574; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_2530 ? _T_2548 : _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2530 | _GEN_38; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2525 ? _T_2529 : _GEN_40; // @[Conditional.scala 40:58]
  reg  bus_cmd_req_hold; // @[el2_ifu_mem_ctl.scala 568:53]
  wire  _T_2590 = ic_act_miss_f | bus_cmd_req_hold; // @[el2_ifu_mem_ctl.scala 564:45]
  reg  ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 565:55]
  wire  _T_2591 = _T_2590 | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 564:64]
  wire  _T_2593 = _T_2591 & _T_2622; // @[el2_ifu_mem_ctl.scala 564:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2595 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 564:133]
  wire  _T_2596 = _T_2595 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 564:164]
  wire  _T_2597 = _T_2596 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 564:184]
  wire  _T_2598 = _T_2597 & miss_pending; // @[el2_ifu_mem_ctl.scala 564:204]
  wire  _T_2599 = ~_T_2598; // @[el2_ifu_mem_ctl.scala 564:112]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 596:45]
  wire  _T_2616 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 599:35]
  wire  _T_2617 = _T_2616 & miss_pending; // @[el2_ifu_mem_ctl.scala 599:53]
  wire  bus_cmd_sent = _T_2617 & _T_2622; // @[el2_ifu_mem_ctl.scala 599:68]
  wire  _T_2602 = ~bus_cmd_sent; // @[el2_ifu_mem_ctl.scala 567:61]
  wire  _T_2603 = _T_2590 & _T_2602; // @[el2_ifu_mem_ctl.scala 567:59]
  wire [2:0] _T_2607 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2609 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2611 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[el2_ifu_mem_ctl.scala 583:57]
  reg  ifu_bus_arvalid_ff; // @[el2_ifu_mem_ctl.scala 585:53]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 597:51]
  wire  _T_2637 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 607:73]
  wire  _T_2638 = _T_2623 & _T_2637; // @[el2_ifu_mem_ctl.scala 607:71]
  wire  _T_2640 = last_data_recieved_ff & _T_1329; // @[el2_ifu_mem_ctl.scala 607:114]
  wire [2:0] _T_2646 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 612:45]
  wire  _T_2650 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 615:48]
  wire  _T_2651 = _T_2650 & miss_pending; // @[el2_ifu_mem_ctl.scala 615:68]
  wire  bus_inc_cmd_beat_cnt = _T_2651 & _T_2622; // @[el2_ifu_mem_ctl.scala 615:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 617:57]
  wire  _T_2655 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 618:31]
  wire  _T_2656 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 618:71]
  wire  _T_2657 = _T_2656 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 618:87]
  wire  _T_2658 = ~_T_2657; // @[el2_ifu_mem_ctl.scala 618:55]
  wire  bus_hold_cmd_beat_cnt = _T_2655 & _T_2658; // @[el2_ifu_mem_ctl.scala 618:53]
  wire  _T_2659 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 619:46]
  wire  bus_cmd_beat_en = _T_2659 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 619:62]
  wire [2:0] _T_2662 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 621:46]
  wire [2:0] _T_2664 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2665 = bus_inc_cmd_beat_cnt ? _T_2662 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2666 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2668 = _T_2664 | _T_2665; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2668 | _T_2666; // @[Mux.scala 27:72]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 633:62]
  wire  _T_2697 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 638:50]
  wire  _T_2698 = io_ifc_dma_access_ok & _T_2697; // @[el2_ifu_mem_ctl.scala 638:47]
  wire  _T_2699 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 638:70]
  wire  _T_2703 = _T_2698 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 639:72]
  wire  _T_2704 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 639:111]
  wire  _T_2705 = _T_2703 & _T_2704; // @[el2_ifu_mem_ctl.scala 639:97]
  wire  ifc_dma_access_q_ok = _T_2705 & _T_2699; // @[el2_ifu_mem_ctl.scala 639:127]
  wire  _T_2708 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 642:40]
  wire  _T_2709 = _T_2708 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 642:58]
  wire  _T_2712 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 643:60]
  wire  _T_2713 = _T_2708 & _T_2712; // @[el2_ifu_mem_ctl.scala 643:58]
  wire  _T_2714 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 643:104]
  wire [2:0] _T_2719 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire  _T_2740 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[33]; // @[el2_lib.scala 259:74]
  wire  _T_2741 = _T_2740 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 259:74]
  wire  _T_2742 = _T_2741 ^ io_dma_mem_wdata[36]; // @[el2_lib.scala 259:74]
  wire  _T_2743 = _T_2742 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 259:74]
  wire  _T_2744 = _T_2743 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 259:74]
  wire  _T_2745 = _T_2744 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2746 = _T_2745 ^ io_dma_mem_wdata[43]; // @[el2_lib.scala 259:74]
  wire  _T_2747 = _T_2746 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 259:74]
  wire  _T_2748 = _T_2747 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 259:74]
  wire  _T_2749 = _T_2748 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2750 = _T_2749 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 259:74]
  wire  _T_2751 = _T_2750 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2752 = _T_2751 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2753 = _T_2752 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2754 = _T_2753 ^ io_dma_mem_wdata[58]; // @[el2_lib.scala 259:74]
  wire  _T_2755 = _T_2754 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 259:74]
  wire  _T_2756 = _T_2755 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 259:74]
  wire  _T_2775 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 259:74]
  wire  _T_2776 = _T_2775 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 259:74]
  wire  _T_2777 = _T_2776 ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 259:74]
  wire  _T_2778 = _T_2777 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 259:74]
  wire  _T_2779 = _T_2778 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 259:74]
  wire  _T_2780 = _T_2779 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2781 = _T_2780 ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 259:74]
  wire  _T_2782 = _T_2781 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 259:74]
  wire  _T_2783 = _T_2782 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 259:74]
  wire  _T_2784 = _T_2783 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2785 = _T_2784 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 259:74]
  wire  _T_2786 = _T_2785 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2787 = _T_2786 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2788 = _T_2787 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2789 = _T_2788 ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 259:74]
  wire  _T_2790 = _T_2789 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 259:74]
  wire  _T_2791 = _T_2790 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 259:74]
  wire  _T_2810 = io_dma_mem_wdata[33] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 259:74]
  wire  _T_2811 = _T_2810 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 259:74]
  wire  _T_2812 = _T_2811 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 259:74]
  wire  _T_2813 = _T_2812 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 259:74]
  wire  _T_2814 = _T_2813 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 259:74]
  wire  _T_2815 = _T_2814 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2816 = _T_2815 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 259:74]
  wire  _T_2817 = _T_2816 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 259:74]
  wire  _T_2818 = _T_2817 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 259:74]
  wire  _T_2819 = _T_2818 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2820 = _T_2819 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 259:74]
  wire  _T_2821 = _T_2820 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2822 = _T_2821 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2823 = _T_2822 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2824 = _T_2823 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 259:74]
  wire  _T_2825 = _T_2824 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 259:74]
  wire  _T_2826 = _T_2825 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 259:74]
  wire  _T_2842 = io_dma_mem_wdata[36] ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 259:74]
  wire  _T_2843 = _T_2842 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 259:74]
  wire  _T_2844 = _T_2843 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 259:74]
  wire  _T_2845 = _T_2844 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 259:74]
  wire  _T_2846 = _T_2845 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 259:74]
  wire  _T_2847 = _T_2846 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 259:74]
  wire  _T_2848 = _T_2847 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 259:74]
  wire  _T_2849 = _T_2848 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 259:74]
  wire  _T_2850 = _T_2849 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 259:74]
  wire  _T_2851 = _T_2850 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2852 = _T_2851 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 259:74]
  wire  _T_2853 = _T_2852 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2854 = _T_2853 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2855 = _T_2854 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2871 = io_dma_mem_wdata[43] ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 259:74]
  wire  _T_2872 = _T_2871 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 259:74]
  wire  _T_2873 = _T_2872 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 259:74]
  wire  _T_2874 = _T_2873 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 259:74]
  wire  _T_2875 = _T_2874 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 259:74]
  wire  _T_2876 = _T_2875 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 259:74]
  wire  _T_2877 = _T_2876 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 259:74]
  wire  _T_2878 = _T_2877 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 259:74]
  wire  _T_2879 = _T_2878 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 259:74]
  wire  _T_2880 = _T_2879 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 259:74]
  wire  _T_2881 = _T_2880 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 259:74]
  wire  _T_2882 = _T_2881 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 259:74]
  wire  _T_2883 = _T_2882 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 259:74]
  wire  _T_2884 = _T_2883 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 259:74]
  wire  _T_2891 = io_dma_mem_wdata[58] ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 259:74]
  wire  _T_2892 = _T_2891 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 259:74]
  wire  _T_2893 = _T_2892 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 259:74]
  wire  _T_2894 = _T_2893 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 259:74]
  wire  _T_2895 = _T_2894 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 259:74]
  wire [5:0] _T_2900 = {_T_2895,_T_2884,_T_2855,_T_2826,_T_2791,_T_2756}; // @[Cat.scala 29:58]
  wire  _T_2901 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 267:13]
  wire  _T_2902 = ^_T_2900; // @[el2_lib.scala 267:23]
  wire  _T_2903 = _T_2901 ^ _T_2902; // @[el2_lib.scala 267:18]
  wire  _T_2924 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[1]; // @[el2_lib.scala 259:74]
  wire  _T_2925 = _T_2924 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 259:74]
  wire  _T_2926 = _T_2925 ^ io_dma_mem_wdata[4]; // @[el2_lib.scala 259:74]
  wire  _T_2927 = _T_2926 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 259:74]
  wire  _T_2928 = _T_2927 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 259:74]
  wire  _T_2929 = _T_2928 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_2930 = _T_2929 ^ io_dma_mem_wdata[11]; // @[el2_lib.scala 259:74]
  wire  _T_2931 = _T_2930 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 259:74]
  wire  _T_2932 = _T_2931 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 259:74]
  wire  _T_2933 = _T_2932 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_2934 = _T_2933 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 259:74]
  wire  _T_2935 = _T_2934 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_2936 = _T_2935 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_2937 = _T_2936 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_2938 = _T_2937 ^ io_dma_mem_wdata[26]; // @[el2_lib.scala 259:74]
  wire  _T_2939 = _T_2938 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 259:74]
  wire  _T_2940 = _T_2939 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 259:74]
  wire  _T_2959 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 259:74]
  wire  _T_2960 = _T_2959 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 259:74]
  wire  _T_2961 = _T_2960 ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 259:74]
  wire  _T_2962 = _T_2961 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 259:74]
  wire  _T_2963 = _T_2962 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 259:74]
  wire  _T_2964 = _T_2963 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_2965 = _T_2964 ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 259:74]
  wire  _T_2966 = _T_2965 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 259:74]
  wire  _T_2967 = _T_2966 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 259:74]
  wire  _T_2968 = _T_2967 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_2969 = _T_2968 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 259:74]
  wire  _T_2970 = _T_2969 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_2971 = _T_2970 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_2972 = _T_2971 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_2973 = _T_2972 ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 259:74]
  wire  _T_2974 = _T_2973 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 259:74]
  wire  _T_2975 = _T_2974 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 259:74]
  wire  _T_2994 = io_dma_mem_wdata[1] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 259:74]
  wire  _T_2995 = _T_2994 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 259:74]
  wire  _T_2996 = _T_2995 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 259:74]
  wire  _T_2997 = _T_2996 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 259:74]
  wire  _T_2998 = _T_2997 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 259:74]
  wire  _T_2999 = _T_2998 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_3000 = _T_2999 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 259:74]
  wire  _T_3001 = _T_3000 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 259:74]
  wire  _T_3002 = _T_3001 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 259:74]
  wire  _T_3003 = _T_3002 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_3004 = _T_3003 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 259:74]
  wire  _T_3005 = _T_3004 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_3006 = _T_3005 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_3007 = _T_3006 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_3008 = _T_3007 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 259:74]
  wire  _T_3009 = _T_3008 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 259:74]
  wire  _T_3010 = _T_3009 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 259:74]
  wire  _T_3026 = io_dma_mem_wdata[4] ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 259:74]
  wire  _T_3027 = _T_3026 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 259:74]
  wire  _T_3028 = _T_3027 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 259:74]
  wire  _T_3029 = _T_3028 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 259:74]
  wire  _T_3030 = _T_3029 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 259:74]
  wire  _T_3031 = _T_3030 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 259:74]
  wire  _T_3032 = _T_3031 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 259:74]
  wire  _T_3033 = _T_3032 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 259:74]
  wire  _T_3034 = _T_3033 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 259:74]
  wire  _T_3035 = _T_3034 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_3036 = _T_3035 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 259:74]
  wire  _T_3037 = _T_3036 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_3038 = _T_3037 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_3039 = _T_3038 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_3055 = io_dma_mem_wdata[11] ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 259:74]
  wire  _T_3056 = _T_3055 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 259:74]
  wire  _T_3057 = _T_3056 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 259:74]
  wire  _T_3058 = _T_3057 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 259:74]
  wire  _T_3059 = _T_3058 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 259:74]
  wire  _T_3060 = _T_3059 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 259:74]
  wire  _T_3061 = _T_3060 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 259:74]
  wire  _T_3062 = _T_3061 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 259:74]
  wire  _T_3063 = _T_3062 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 259:74]
  wire  _T_3064 = _T_3063 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 259:74]
  wire  _T_3065 = _T_3064 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 259:74]
  wire  _T_3066 = _T_3065 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 259:74]
  wire  _T_3067 = _T_3066 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 259:74]
  wire  _T_3068 = _T_3067 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 259:74]
  wire  _T_3075 = io_dma_mem_wdata[26] ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 259:74]
  wire  _T_3076 = _T_3075 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 259:74]
  wire  _T_3077 = _T_3076 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 259:74]
  wire  _T_3078 = _T_3077 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 259:74]
  wire  _T_3079 = _T_3078 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 259:74]
  wire [5:0] _T_3084 = {_T_3079,_T_3068,_T_3039,_T_3010,_T_2975,_T_2940}; // @[Cat.scala 29:58]
  wire  _T_3085 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 267:13]
  wire  _T_3086 = ^_T_3084; // @[el2_lib.scala 267:23]
  wire  _T_3087 = _T_3085 ^ _T_3086; // @[el2_lib.scala 267:18]
  wire [6:0] _T_3088 = {_T_3087,_T_3079,_T_3068,_T_3039,_T_3010,_T_2975,_T_2940}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2903,_T_2895,_T_2884,_T_2855,_T_2826,_T_2791,_T_2756,_T_3088}; // @[Cat.scala 29:58]
  wire  _T_3090 = ~_T_2708; // @[el2_ifu_mem_ctl.scala 649:45]
  wire  _T_3091 = iccm_correct_ecc & _T_3090; // @[el2_ifu_mem_ctl.scala 649:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3092 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3099 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 663:53]
  wire  _T_3434 = _T_3346[5:0] == 6'h27; // @[el2_lib.scala 339:41]
  wire  _T_3432 = _T_3346[5:0] == 6'h26; // @[el2_lib.scala 339:41]
  wire  _T_3430 = _T_3346[5:0] == 6'h25; // @[el2_lib.scala 339:41]
  wire  _T_3428 = _T_3346[5:0] == 6'h24; // @[el2_lib.scala 339:41]
  wire  _T_3426 = _T_3346[5:0] == 6'h23; // @[el2_lib.scala 339:41]
  wire  _T_3424 = _T_3346[5:0] == 6'h22; // @[el2_lib.scala 339:41]
  wire  _T_3422 = _T_3346[5:0] == 6'h21; // @[el2_lib.scala 339:41]
  wire  _T_3420 = _T_3346[5:0] == 6'h20; // @[el2_lib.scala 339:41]
  wire  _T_3418 = _T_3346[5:0] == 6'h1f; // @[el2_lib.scala 339:41]
  wire  _T_3416 = _T_3346[5:0] == 6'h1e; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3492 = {_T_3434,_T_3432,_T_3430,_T_3428,_T_3426,_T_3424,_T_3422,_T_3420,_T_3418,_T_3416}; // @[el2_lib.scala 342:69]
  wire  _T_3414 = _T_3346[5:0] == 6'h1d; // @[el2_lib.scala 339:41]
  wire  _T_3412 = _T_3346[5:0] == 6'h1c; // @[el2_lib.scala 339:41]
  wire  _T_3410 = _T_3346[5:0] == 6'h1b; // @[el2_lib.scala 339:41]
  wire  _T_3408 = _T_3346[5:0] == 6'h1a; // @[el2_lib.scala 339:41]
  wire  _T_3406 = _T_3346[5:0] == 6'h19; // @[el2_lib.scala 339:41]
  wire  _T_3404 = _T_3346[5:0] == 6'h18; // @[el2_lib.scala 339:41]
  wire  _T_3402 = _T_3346[5:0] == 6'h17; // @[el2_lib.scala 339:41]
  wire  _T_3400 = _T_3346[5:0] == 6'h16; // @[el2_lib.scala 339:41]
  wire  _T_3398 = _T_3346[5:0] == 6'h15; // @[el2_lib.scala 339:41]
  wire  _T_3396 = _T_3346[5:0] == 6'h14; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3483 = {_T_3414,_T_3412,_T_3410,_T_3408,_T_3406,_T_3404,_T_3402,_T_3400,_T_3398,_T_3396}; // @[el2_lib.scala 342:69]
  wire  _T_3394 = _T_3346[5:0] == 6'h13; // @[el2_lib.scala 339:41]
  wire  _T_3392 = _T_3346[5:0] == 6'h12; // @[el2_lib.scala 339:41]
  wire  _T_3390 = _T_3346[5:0] == 6'h11; // @[el2_lib.scala 339:41]
  wire  _T_3388 = _T_3346[5:0] == 6'h10; // @[el2_lib.scala 339:41]
  wire  _T_3386 = _T_3346[5:0] == 6'hf; // @[el2_lib.scala 339:41]
  wire  _T_3384 = _T_3346[5:0] == 6'he; // @[el2_lib.scala 339:41]
  wire  _T_3382 = _T_3346[5:0] == 6'hd; // @[el2_lib.scala 339:41]
  wire  _T_3380 = _T_3346[5:0] == 6'hc; // @[el2_lib.scala 339:41]
  wire  _T_3378 = _T_3346[5:0] == 6'hb; // @[el2_lib.scala 339:41]
  wire  _T_3376 = _T_3346[5:0] == 6'ha; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3473 = {_T_3394,_T_3392,_T_3390,_T_3388,_T_3386,_T_3384,_T_3382,_T_3380,_T_3378,_T_3376}; // @[el2_lib.scala 342:69]
  wire  _T_3374 = _T_3346[5:0] == 6'h9; // @[el2_lib.scala 339:41]
  wire  _T_3372 = _T_3346[5:0] == 6'h8; // @[el2_lib.scala 339:41]
  wire  _T_3370 = _T_3346[5:0] == 6'h7; // @[el2_lib.scala 339:41]
  wire  _T_3368 = _T_3346[5:0] == 6'h6; // @[el2_lib.scala 339:41]
  wire  _T_3366 = _T_3346[5:0] == 6'h5; // @[el2_lib.scala 339:41]
  wire  _T_3364 = _T_3346[5:0] == 6'h4; // @[el2_lib.scala 339:41]
  wire  _T_3362 = _T_3346[5:0] == 6'h3; // @[el2_lib.scala 339:41]
  wire  _T_3360 = _T_3346[5:0] == 6'h2; // @[el2_lib.scala 339:41]
  wire  _T_3358 = _T_3346[5:0] == 6'h1; // @[el2_lib.scala 339:41]
  wire [18:0] _T_3474 = {_T_3473,_T_3374,_T_3372,_T_3370,_T_3368,_T_3366,_T_3364,_T_3362,_T_3360,_T_3358}; // @[el2_lib.scala 342:69]
  wire [38:0] _T_3494 = {_T_3492,_T_3483,_T_3474}; // @[el2_lib.scala 342:69]
  wire [7:0] _T_3449 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3455 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3449}; // @[Cat.scala 29:58]
  wire [38:0] _T_3495 = _T_3494 ^ _T_3455; // @[el2_lib.scala 342:76]
  wire [38:0] _T_3496 = _T_3350 ? _T_3495 : _T_3455; // @[el2_lib.scala 342:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3496[37:32],_T_3496[30:16],_T_3496[14:8],_T_3496[6:4],_T_3496[2]}; // @[Cat.scala 29:58]
  wire  _T_3819 = _T_3731[5:0] == 6'h27; // @[el2_lib.scala 339:41]
  wire  _T_3817 = _T_3731[5:0] == 6'h26; // @[el2_lib.scala 339:41]
  wire  _T_3815 = _T_3731[5:0] == 6'h25; // @[el2_lib.scala 339:41]
  wire  _T_3813 = _T_3731[5:0] == 6'h24; // @[el2_lib.scala 339:41]
  wire  _T_3811 = _T_3731[5:0] == 6'h23; // @[el2_lib.scala 339:41]
  wire  _T_3809 = _T_3731[5:0] == 6'h22; // @[el2_lib.scala 339:41]
  wire  _T_3807 = _T_3731[5:0] == 6'h21; // @[el2_lib.scala 339:41]
  wire  _T_3805 = _T_3731[5:0] == 6'h20; // @[el2_lib.scala 339:41]
  wire  _T_3803 = _T_3731[5:0] == 6'h1f; // @[el2_lib.scala 339:41]
  wire  _T_3801 = _T_3731[5:0] == 6'h1e; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3877 = {_T_3819,_T_3817,_T_3815,_T_3813,_T_3811,_T_3809,_T_3807,_T_3805,_T_3803,_T_3801}; // @[el2_lib.scala 342:69]
  wire  _T_3799 = _T_3731[5:0] == 6'h1d; // @[el2_lib.scala 339:41]
  wire  _T_3797 = _T_3731[5:0] == 6'h1c; // @[el2_lib.scala 339:41]
  wire  _T_3795 = _T_3731[5:0] == 6'h1b; // @[el2_lib.scala 339:41]
  wire  _T_3793 = _T_3731[5:0] == 6'h1a; // @[el2_lib.scala 339:41]
  wire  _T_3791 = _T_3731[5:0] == 6'h19; // @[el2_lib.scala 339:41]
  wire  _T_3789 = _T_3731[5:0] == 6'h18; // @[el2_lib.scala 339:41]
  wire  _T_3787 = _T_3731[5:0] == 6'h17; // @[el2_lib.scala 339:41]
  wire  _T_3785 = _T_3731[5:0] == 6'h16; // @[el2_lib.scala 339:41]
  wire  _T_3783 = _T_3731[5:0] == 6'h15; // @[el2_lib.scala 339:41]
  wire  _T_3781 = _T_3731[5:0] == 6'h14; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3868 = {_T_3799,_T_3797,_T_3795,_T_3793,_T_3791,_T_3789,_T_3787,_T_3785,_T_3783,_T_3781}; // @[el2_lib.scala 342:69]
  wire  _T_3779 = _T_3731[5:0] == 6'h13; // @[el2_lib.scala 339:41]
  wire  _T_3777 = _T_3731[5:0] == 6'h12; // @[el2_lib.scala 339:41]
  wire  _T_3775 = _T_3731[5:0] == 6'h11; // @[el2_lib.scala 339:41]
  wire  _T_3773 = _T_3731[5:0] == 6'h10; // @[el2_lib.scala 339:41]
  wire  _T_3771 = _T_3731[5:0] == 6'hf; // @[el2_lib.scala 339:41]
  wire  _T_3769 = _T_3731[5:0] == 6'he; // @[el2_lib.scala 339:41]
  wire  _T_3767 = _T_3731[5:0] == 6'hd; // @[el2_lib.scala 339:41]
  wire  _T_3765 = _T_3731[5:0] == 6'hc; // @[el2_lib.scala 339:41]
  wire  _T_3763 = _T_3731[5:0] == 6'hb; // @[el2_lib.scala 339:41]
  wire  _T_3761 = _T_3731[5:0] == 6'ha; // @[el2_lib.scala 339:41]
  wire [9:0] _T_3858 = {_T_3779,_T_3777,_T_3775,_T_3773,_T_3771,_T_3769,_T_3767,_T_3765,_T_3763,_T_3761}; // @[el2_lib.scala 342:69]
  wire  _T_3759 = _T_3731[5:0] == 6'h9; // @[el2_lib.scala 339:41]
  wire  _T_3757 = _T_3731[5:0] == 6'h8; // @[el2_lib.scala 339:41]
  wire  _T_3755 = _T_3731[5:0] == 6'h7; // @[el2_lib.scala 339:41]
  wire  _T_3753 = _T_3731[5:0] == 6'h6; // @[el2_lib.scala 339:41]
  wire  _T_3751 = _T_3731[5:0] == 6'h5; // @[el2_lib.scala 339:41]
  wire  _T_3749 = _T_3731[5:0] == 6'h4; // @[el2_lib.scala 339:41]
  wire  _T_3747 = _T_3731[5:0] == 6'h3; // @[el2_lib.scala 339:41]
  wire  _T_3745 = _T_3731[5:0] == 6'h2; // @[el2_lib.scala 339:41]
  wire  _T_3743 = _T_3731[5:0] == 6'h1; // @[el2_lib.scala 339:41]
  wire [18:0] _T_3859 = {_T_3858,_T_3759,_T_3757,_T_3755,_T_3753,_T_3751,_T_3749,_T_3747,_T_3745,_T_3743}; // @[el2_lib.scala 342:69]
  wire [38:0] _T_3879 = {_T_3877,_T_3868,_T_3859}; // @[el2_lib.scala 342:69]
  wire [7:0] _T_3834 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3840 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3834}; // @[Cat.scala 29:58]
  wire [38:0] _T_3880 = _T_3879 ^ _T_3840; // @[el2_lib.scala 342:76]
  wire [38:0] _T_3881 = _T_3735 ? _T_3880 : _T_3840; // @[el2_lib.scala 342:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3881[37:32],_T_3881[30:16],_T_3881[14:8],_T_3881[6:4],_T_3881[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 655:35]
  wire  _T_3354 = ~_T_3346[6]; // @[el2_lib.scala 335:55]
  wire  _T_3355 = _T_3348 & _T_3354; // @[el2_lib.scala 335:53]
  wire  _T_3739 = ~_T_3731[6]; // @[el2_lib.scala 335:55]
  wire  _T_3740 = _T_3733 & _T_3739; // @[el2_lib.scala 335:53]
  wire [1:0] iccm_double_ecc_error = {_T_3355,_T_3740}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 657:53]
  wire [63:0] _T_3103 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3104 = {iccm_dma_rdata_1_muxed,_T_3496[37:32],_T_3496[30:16],_T_3496[14:8],_T_3496[6:4],_T_3496[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 659:54]
  reg [2:0] iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 660:74]
  reg  iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 665:76]
  reg  iccm_dma_ecc_error; // @[el2_ifu_mem_ctl.scala 667:74]
  reg [63:0] iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 669:75]
  wire  _T_3109 = _T_2708 & _T_2697; // @[el2_ifu_mem_ctl.scala 672:65]
  wire  _T_3113 = _T_3090 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 673:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3114 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [14:0] _T_3116 = _T_3113 ? _T_3114 : io_ifc_fetch_addr_bf[14:0]; // @[el2_ifu_mem_ctl.scala 673:8]
  wire  _T_3508 = _T_3346 == 7'h40; // @[el2_lib.scala 345:62]
  wire  _T_3509 = _T_3496[38] ^ _T_3508; // @[el2_lib.scala 345:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3509,_T_3496[31],_T_3496[15],_T_3496[7],_T_3496[3],_T_3496[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3893 = _T_3731 == 7'h40; // @[el2_lib.scala 345:62]
  wire  _T_3894 = _T_3881[38] ^ _T_3893; // @[el2_lib.scala 345:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3894,_T_3881[31],_T_3881[15],_T_3881[7],_T_3881[3],_T_3881[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3910 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 685:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 687:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 688:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 696:62]
  wire  _T_3918 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 690:76]
  wire  _T_3919 = io_iccm_rd_ecc_single_err & _T_3918; // @[el2_ifu_mem_ctl.scala 690:74]
  wire  _T_3921 = _T_3919 & _T_319; // @[el2_ifu_mem_ctl.scala 690:104]
  wire  iccm_ecc_write_status = _T_3921 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 690:127]
  wire  _T_3922 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 691:67]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 695:51]
  wire [13:0] _T_3927 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 694:102]
  wire [38:0] _T_3931 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3936 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 699:41]
  wire  _T_3937 = io_ifc_fetch_req_bf & _T_3936; // @[el2_ifu_mem_ctl.scala 699:39]
  wire  _T_3938 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 699:72]
  wire  _T_3939 = _T_3937 & _T_3938; // @[el2_ifu_mem_ctl.scala 699:70]
  wire  _T_3941 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 700:34]
  wire  _T_3942 = _T_2267 & _T_3941; // @[el2_ifu_mem_ctl.scala 700:32]
  wire  _T_3945 = _T_2283 & _T_3941; // @[el2_ifu_mem_ctl.scala 701:37]
  wire  _T_3946 = _T_3942 | _T_3945; // @[el2_ifu_mem_ctl.scala 700:88]
  wire  _T_3947 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 702:19]
  wire  _T_3949 = _T_3947 & _T_3941; // @[el2_ifu_mem_ctl.scala 702:41]
  wire  _T_3950 = _T_3946 | _T_3949; // @[el2_ifu_mem_ctl.scala 701:88]
  wire  _T_3951 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 703:19]
  wire  _T_3953 = _T_3951 & _T_3941; // @[el2_ifu_mem_ctl.scala 703:35]
  wire  _T_3954 = _T_3950 | _T_3953; // @[el2_ifu_mem_ctl.scala 702:88]
  wire  _T_3957 = _T_2282 & _T_3941; // @[el2_ifu_mem_ctl.scala 704:38]
  wire  _T_3958 = _T_3954 | _T_3957; // @[el2_ifu_mem_ctl.scala 703:88]
  wire  _T_3960 = _T_2283 & miss_state_en; // @[el2_ifu_mem_ctl.scala 705:37]
  wire  _T_3961 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 705:71]
  wire  _T_3962 = _T_3960 & _T_3961; // @[el2_ifu_mem_ctl.scala 705:54]
  wire  _T_3963 = _T_3958 | _T_3962; // @[el2_ifu_mem_ctl.scala 704:57]
  wire  _T_3964 = ~_T_3963; // @[el2_ifu_mem_ctl.scala 700:5]
  wire  _T_3965 = _T_3939 & _T_3964; // @[el2_ifu_mem_ctl.scala 699:96]
  wire  _T_3966 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 706:28]
  wire  _T_3968 = _T_3966 & _T_3936; // @[el2_ifu_mem_ctl.scala 706:50]
  wire  _T_3970 = _T_3968 & _T_3938; // @[el2_ifu_mem_ctl.scala 706:81]
  wire [1:0] _T_3973 = write_ic_16_bytes ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9779 = bus_ifu_wr_en_ff_q & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 801:74]
  wire  bus_wren_1 = _T_9779 & miss_pending; // @[el2_ifu_mem_ctl.scala 801:98]
  wire  _T_9778 = bus_ifu_wr_en_ff_q & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 801:74]
  wire  bus_wren_0 = _T_9778 & miss_pending; // @[el2_ifu_mem_ctl.scala 801:98]
  wire [1:0] bus_ic_wr_en = {bus_wren_1,bus_wren_0}; // @[Cat.scala 29:58]
  wire  _T_3979 = ~_T_108; // @[el2_ifu_mem_ctl.scala 709:106]
  wire  _T_3980 = _T_2267 & _T_3979; // @[el2_ifu_mem_ctl.scala 709:104]
  wire  _T_3981 = _T_2283 | _T_3980; // @[el2_ifu_mem_ctl.scala 709:77]
  wire  _T_3985 = ~_T_51; // @[el2_ifu_mem_ctl.scala 709:172]
  wire  _T_3986 = _T_3981 & _T_3985; // @[el2_ifu_mem_ctl.scala 709:170]
  wire  _T_3987 = ~_T_3986; // @[el2_ifu_mem_ctl.scala 709:44]
  wire  _T_3991 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 712:64]
  wire  _T_3992 = ~_T_3991; // @[el2_ifu_mem_ctl.scala 712:50]
  wire  _T_3993 = _T_276 & _T_3992; // @[el2_ifu_mem_ctl.scala 712:48]
  wire  _T_3994 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 712:81]
  wire  ic_valid = _T_3993 & _T_3994; // @[el2_ifu_mem_ctl.scala 712:79]
  wire  _T_3996 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 713:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 716:14]
  wire  _T_3999 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 719:74]
  wire  _T_9776 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 800:45]
  wire  way_status_wr_en = _T_9776 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 800:58]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 721:14]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 796:41]
  reg  way_status_new_ff; // @[el2_ifu_mem_ctl.scala 727:14]
  wire  _T_4019 = ifu_status_wr_addr_ff[2:0] == 3'h0; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4020 = _T_4019 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 733:136]
  wire  _T_4023 = ifu_status_wr_addr_ff[2:0] == 3'h1; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4024 = _T_4023 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 733:136]
  wire  _T_4027 = ifu_status_wr_addr_ff[2:0] == 3'h2; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4028 = _T_4027 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 733:136]
  wire  _T_4031 = ifu_status_wr_addr_ff[2:0] == 3'h3; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4032 = _T_4031 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 733:136]
  wire  _T_4035 = ifu_status_wr_addr_ff[2:0] == 3'h4; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4036 = _T_4035 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 733:136]
  wire  _T_4039 = ifu_status_wr_addr_ff[2:0] == 3'h5; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4040 = _T_4039 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 733:136]
  wire  _T_4043 = ifu_status_wr_addr_ff[2:0] == 3'h6; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4044 = _T_4043 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 733:136]
  wire  _T_4047 = ifu_status_wr_addr_ff[2:0] == 3'h7; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4048 = _T_4047 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 733:136]
  wire  _T_9782 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 803:84]
  wire  _T_9783 = _T_9782 & miss_pending; // @[el2_ifu_mem_ctl.scala 803:108]
  wire  bus_wren_last_1 = _T_9783 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 803:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 804:84]
  wire  _T_9785 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 805:73]
  wire  _T_9780 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 803:84]
  wire  _T_9781 = _T_9780 & miss_pending; // @[el2_ifu_mem_ctl.scala 803:108]
  wire  bus_wren_last_0 = _T_9781 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 803:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 804:84]
  wire  _T_9784 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 805:73]
  wire [1:0] ifu_tag_wren = {_T_9785,_T_9784}; // @[Cat.scala 29:58]
  wire [1:0] _T_9820 = _T_3999 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_9820 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 839:90]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 748:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 752:14]
  wire  _T_5062 = ifu_ic_rw_int_addr_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 756:78]
  wire  _T_5064 = _T_5062 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 756:87]
  wire  _T_5066 = perr_ic_index_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 757:70]
  wire  _T_5068 = _T_5066 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:79]
  wire  _T_5069 = _T_5064 | _T_5068; // @[el2_ifu_mem_ctl.scala 756:109]
  wire  _T_5070 = _T_5069 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5074 = _T_5062 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 756:87]
  wire  _T_5078 = _T_5066 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:79]
  wire  _T_5079 = _T_5074 | _T_5078; // @[el2_ifu_mem_ctl.scala 756:109]
  wire  _T_5080 = _T_5079 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:102]
  wire [1:0] tag_valid_clken_0 = {_T_5080,_T_5070}; // @[Cat.scala 29:58]
  wire  _T_5082 = ifu_ic_rw_int_addr_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 756:78]
  wire  _T_5084 = _T_5082 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 756:87]
  wire  _T_5086 = perr_ic_index_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 757:70]
  wire  _T_5088 = _T_5086 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:79]
  wire  _T_5089 = _T_5084 | _T_5088; // @[el2_ifu_mem_ctl.scala 756:109]
  wire  _T_5090 = _T_5089 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5094 = _T_5082 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 756:87]
  wire  _T_5098 = _T_5086 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:79]
  wire  _T_5099 = _T_5094 | _T_5098; // @[el2_ifu_mem_ctl.scala 756:109]
  wire  _T_5100 = _T_5099 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:102]
  wire [1:0] tag_valid_clken_1 = {_T_5100,_T_5090}; // @[Cat.scala 29:58]
  wire  _T_5102 = ifu_ic_rw_int_addr_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 756:78]
  wire  _T_5104 = _T_5102 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 756:87]
  wire  _T_5106 = perr_ic_index_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 757:70]
  wire  _T_5108 = _T_5106 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:79]
  wire  _T_5109 = _T_5104 | _T_5108; // @[el2_ifu_mem_ctl.scala 756:109]
  wire  _T_5110 = _T_5109 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5114 = _T_5102 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 756:87]
  wire  _T_5118 = _T_5106 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:79]
  wire  _T_5119 = _T_5114 | _T_5118; // @[el2_ifu_mem_ctl.scala 756:109]
  wire  _T_5120 = _T_5119 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:102]
  wire [1:0] tag_valid_clken_2 = {_T_5120,_T_5110}; // @[Cat.scala 29:58]
  wire  _T_5122 = ifu_ic_rw_int_addr_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 756:78]
  wire  _T_5124 = _T_5122 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 756:87]
  wire  _T_5126 = perr_ic_index_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 757:70]
  wire  _T_5128 = _T_5126 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:79]
  wire  _T_5129 = _T_5124 | _T_5128; // @[el2_ifu_mem_ctl.scala 756:109]
  wire  _T_5130 = _T_5129 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5134 = _T_5122 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 756:87]
  wire  _T_5138 = _T_5126 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:79]
  wire  _T_5139 = _T_5134 | _T_5138; // @[el2_ifu_mem_ctl.scala 756:109]
  wire  _T_5140 = _T_5139 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:102]
  wire [1:0] tag_valid_clken_3 = {_T_5140,_T_5130}; // @[Cat.scala 29:58]
  wire  _T_5151 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 765:97]
  wire  _T_5152 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 765:124]
  wire  _T_5153 = _T_5151 & _T_5152; // @[el2_ifu_mem_ctl.scala 765:122]
  wire  _T_5156 = _T_4670 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5157 = perr_ic_index_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5159 = _T_5157 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5160 = _T_5156 | _T_5159; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5161 = _T_5160 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5171 = _T_4671 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5172 = perr_ic_index_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5174 = _T_5172 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5175 = _T_5171 | _T_5174; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5176 = _T_5175 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5186 = _T_4672 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5187 = perr_ic_index_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5189 = _T_5187 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5190 = _T_5186 | _T_5189; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5191 = _T_5190 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5201 = _T_4673 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5202 = perr_ic_index_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5204 = _T_5202 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5205 = _T_5201 | _T_5204; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5206 = _T_5205 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5216 = _T_4674 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5217 = perr_ic_index_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5219 = _T_5217 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5220 = _T_5216 | _T_5219; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5221 = _T_5220 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5231 = _T_4675 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5232 = perr_ic_index_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5234 = _T_5232 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5235 = _T_5231 | _T_5234; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5236 = _T_5235 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5246 = _T_4676 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5247 = perr_ic_index_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5249 = _T_5247 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5250 = _T_5246 | _T_5249; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5251 = _T_5250 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5261 = _T_4677 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5262 = perr_ic_index_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5264 = _T_5262 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5265 = _T_5261 | _T_5264; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5266 = _T_5265 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5276 = _T_4678 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5277 = perr_ic_index_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5279 = _T_5277 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5280 = _T_5276 | _T_5279; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5281 = _T_5280 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5291 = _T_4679 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5292 = perr_ic_index_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5294 = _T_5292 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5295 = _T_5291 | _T_5294; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5296 = _T_5295 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5306 = _T_4680 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5307 = perr_ic_index_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5309 = _T_5307 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5310 = _T_5306 | _T_5309; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5311 = _T_5310 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5321 = _T_4681 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5322 = perr_ic_index_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5324 = _T_5322 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5325 = _T_5321 | _T_5324; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5326 = _T_5325 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5336 = _T_4682 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5337 = perr_ic_index_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5339 = _T_5337 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5340 = _T_5336 | _T_5339; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5341 = _T_5340 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5351 = _T_4683 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5352 = perr_ic_index_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5354 = _T_5352 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5355 = _T_5351 | _T_5354; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5356 = _T_5355 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5366 = _T_4684 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5367 = perr_ic_index_ff == 7'he; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5369 = _T_5367 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5370 = _T_5366 | _T_5369; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5371 = _T_5370 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5381 = _T_4685 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5382 = perr_ic_index_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5384 = _T_5382 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5385 = _T_5381 | _T_5384; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5386 = _T_5385 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5396 = _T_4686 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5397 = perr_ic_index_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5399 = _T_5397 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5400 = _T_5396 | _T_5399; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5401 = _T_5400 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5411 = _T_4687 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5412 = perr_ic_index_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5414 = _T_5412 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5415 = _T_5411 | _T_5414; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5416 = _T_5415 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5426 = _T_4688 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5427 = perr_ic_index_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5429 = _T_5427 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5430 = _T_5426 | _T_5429; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5431 = _T_5430 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5441 = _T_4689 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5442 = perr_ic_index_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5444 = _T_5442 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5445 = _T_5441 | _T_5444; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5446 = _T_5445 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5456 = _T_4690 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5457 = perr_ic_index_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5459 = _T_5457 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5460 = _T_5456 | _T_5459; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5461 = _T_5460 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5471 = _T_4691 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5472 = perr_ic_index_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5474 = _T_5472 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5475 = _T_5471 | _T_5474; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5476 = _T_5475 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5486 = _T_4692 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5487 = perr_ic_index_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5489 = _T_5487 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5490 = _T_5486 | _T_5489; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5491 = _T_5490 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5501 = _T_4693 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5502 = perr_ic_index_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5504 = _T_5502 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5505 = _T_5501 | _T_5504; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5506 = _T_5505 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5516 = _T_4694 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5517 = perr_ic_index_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5519 = _T_5517 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5520 = _T_5516 | _T_5519; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5521 = _T_5520 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5531 = _T_4695 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5532 = perr_ic_index_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5534 = _T_5532 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5535 = _T_5531 | _T_5534; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5536 = _T_5535 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5546 = _T_4696 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5547 = perr_ic_index_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5549 = _T_5547 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5550 = _T_5546 | _T_5549; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5551 = _T_5550 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5561 = _T_4697 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5562 = perr_ic_index_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5564 = _T_5562 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5565 = _T_5561 | _T_5564; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5566 = _T_5565 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5576 = _T_4698 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5577 = perr_ic_index_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5579 = _T_5577 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5580 = _T_5576 | _T_5579; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5581 = _T_5580 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5591 = _T_4699 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5592 = perr_ic_index_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5594 = _T_5592 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5595 = _T_5591 | _T_5594; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5596 = _T_5595 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5606 = _T_4700 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5607 = perr_ic_index_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5609 = _T_5607 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5610 = _T_5606 | _T_5609; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5611 = _T_5610 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5621 = _T_4701 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5622 = perr_ic_index_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_5624 = _T_5622 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5625 = _T_5621 | _T_5624; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5626 = _T_5625 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5636 = _T_4670 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5639 = _T_5157 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5640 = _T_5636 | _T_5639; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5641 = _T_5640 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5651 = _T_4671 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5654 = _T_5172 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5655 = _T_5651 | _T_5654; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5656 = _T_5655 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5666 = _T_4672 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5669 = _T_5187 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5670 = _T_5666 | _T_5669; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5671 = _T_5670 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5681 = _T_4673 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5684 = _T_5202 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5685 = _T_5681 | _T_5684; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5686 = _T_5685 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5696 = _T_4674 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5699 = _T_5217 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5700 = _T_5696 | _T_5699; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5701 = _T_5700 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5711 = _T_4675 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5714 = _T_5232 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5715 = _T_5711 | _T_5714; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5716 = _T_5715 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5726 = _T_4676 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5729 = _T_5247 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5730 = _T_5726 | _T_5729; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5731 = _T_5730 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5741 = _T_4677 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5744 = _T_5262 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5745 = _T_5741 | _T_5744; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5746 = _T_5745 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5756 = _T_4678 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5759 = _T_5277 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5760 = _T_5756 | _T_5759; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5761 = _T_5760 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5771 = _T_4679 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5774 = _T_5292 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5775 = _T_5771 | _T_5774; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5776 = _T_5775 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5786 = _T_4680 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5789 = _T_5307 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5790 = _T_5786 | _T_5789; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5791 = _T_5790 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5801 = _T_4681 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5804 = _T_5322 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5805 = _T_5801 | _T_5804; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5806 = _T_5805 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5816 = _T_4682 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5819 = _T_5337 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5820 = _T_5816 | _T_5819; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5821 = _T_5820 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5831 = _T_4683 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5834 = _T_5352 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5835 = _T_5831 | _T_5834; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5836 = _T_5835 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5846 = _T_4684 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5849 = _T_5367 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5850 = _T_5846 | _T_5849; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5851 = _T_5850 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5861 = _T_4685 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5864 = _T_5382 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5865 = _T_5861 | _T_5864; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5866 = _T_5865 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5876 = _T_4686 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5879 = _T_5397 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5880 = _T_5876 | _T_5879; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5881 = _T_5880 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5891 = _T_4687 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5894 = _T_5412 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5895 = _T_5891 | _T_5894; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5896 = _T_5895 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5906 = _T_4688 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5909 = _T_5427 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5910 = _T_5906 | _T_5909; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5911 = _T_5910 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5921 = _T_4689 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5924 = _T_5442 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5925 = _T_5921 | _T_5924; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5926 = _T_5925 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5936 = _T_4690 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5939 = _T_5457 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5940 = _T_5936 | _T_5939; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5941 = _T_5940 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5951 = _T_4691 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5954 = _T_5472 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5955 = _T_5951 | _T_5954; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5956 = _T_5955 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5966 = _T_4692 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5969 = _T_5487 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5970 = _T_5966 | _T_5969; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5971 = _T_5970 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5981 = _T_4693 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5984 = _T_5502 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_5985 = _T_5981 | _T_5984; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_5986 = _T_5985 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_5996 = _T_4694 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_5999 = _T_5517 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6000 = _T_5996 | _T_5999; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6001 = _T_6000 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6011 = _T_4695 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6014 = _T_5532 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6015 = _T_6011 | _T_6014; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6016 = _T_6015 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6026 = _T_4696 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6029 = _T_5547 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6030 = _T_6026 | _T_6029; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6031 = _T_6030 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6041 = _T_4697 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6044 = _T_5562 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6045 = _T_6041 | _T_6044; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6046 = _T_6045 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6056 = _T_4698 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6059 = _T_5577 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6060 = _T_6056 | _T_6059; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6061 = _T_6060 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6071 = _T_4699 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6074 = _T_5592 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6075 = _T_6071 | _T_6074; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6076 = _T_6075 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6086 = _T_4700 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6089 = _T_5607 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6090 = _T_6086 | _T_6089; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6091 = _T_6090 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6101 = _T_4701 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6104 = _T_5622 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6105 = _T_6101 | _T_6104; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6106 = _T_6105 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6116 = _T_4702 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6117 = perr_ic_index_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6119 = _T_6117 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6120 = _T_6116 | _T_6119; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6121 = _T_6120 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6131 = _T_4703 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6132 = perr_ic_index_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6134 = _T_6132 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6135 = _T_6131 | _T_6134; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6136 = _T_6135 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6146 = _T_4704 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6147 = perr_ic_index_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6149 = _T_6147 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6150 = _T_6146 | _T_6149; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6151 = _T_6150 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6161 = _T_4705 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6162 = perr_ic_index_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6164 = _T_6162 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6165 = _T_6161 | _T_6164; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6166 = _T_6165 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6176 = _T_4706 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6177 = perr_ic_index_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6179 = _T_6177 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6180 = _T_6176 | _T_6179; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6181 = _T_6180 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6191 = _T_4707 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6192 = perr_ic_index_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6194 = _T_6192 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6195 = _T_6191 | _T_6194; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6196 = _T_6195 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6206 = _T_4708 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6207 = perr_ic_index_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6209 = _T_6207 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6210 = _T_6206 | _T_6209; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6211 = _T_6210 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6221 = _T_4709 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6222 = perr_ic_index_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6224 = _T_6222 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6225 = _T_6221 | _T_6224; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6226 = _T_6225 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6236 = _T_4710 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6237 = perr_ic_index_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6239 = _T_6237 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6240 = _T_6236 | _T_6239; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6241 = _T_6240 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6251 = _T_4711 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6252 = perr_ic_index_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6254 = _T_6252 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6255 = _T_6251 | _T_6254; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6256 = _T_6255 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6266 = _T_4712 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6267 = perr_ic_index_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6269 = _T_6267 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6270 = _T_6266 | _T_6269; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6271 = _T_6270 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6281 = _T_4713 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6282 = perr_ic_index_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6284 = _T_6282 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6285 = _T_6281 | _T_6284; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6286 = _T_6285 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6296 = _T_4714 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6297 = perr_ic_index_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6299 = _T_6297 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6300 = _T_6296 | _T_6299; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6301 = _T_6300 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6311 = _T_4715 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6312 = perr_ic_index_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6314 = _T_6312 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6315 = _T_6311 | _T_6314; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6316 = _T_6315 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6326 = _T_4716 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6327 = perr_ic_index_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6329 = _T_6327 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6330 = _T_6326 | _T_6329; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6331 = _T_6330 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6341 = _T_4717 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6342 = perr_ic_index_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6344 = _T_6342 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6345 = _T_6341 | _T_6344; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6346 = _T_6345 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6356 = _T_4718 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6357 = perr_ic_index_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6359 = _T_6357 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6360 = _T_6356 | _T_6359; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6361 = _T_6360 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6371 = _T_4719 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6372 = perr_ic_index_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6374 = _T_6372 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6375 = _T_6371 | _T_6374; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6376 = _T_6375 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6386 = _T_4720 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6387 = perr_ic_index_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6389 = _T_6387 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6390 = _T_6386 | _T_6389; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6391 = _T_6390 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6401 = _T_4721 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6402 = perr_ic_index_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6404 = _T_6402 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6405 = _T_6401 | _T_6404; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6406 = _T_6405 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6416 = _T_4722 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6417 = perr_ic_index_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6419 = _T_6417 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6420 = _T_6416 | _T_6419; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6421 = _T_6420 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6431 = _T_4723 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6432 = perr_ic_index_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6434 = _T_6432 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6435 = _T_6431 | _T_6434; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6436 = _T_6435 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6446 = _T_4724 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6447 = perr_ic_index_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6449 = _T_6447 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6450 = _T_6446 | _T_6449; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6451 = _T_6450 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6461 = _T_4725 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6462 = perr_ic_index_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6464 = _T_6462 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6465 = _T_6461 | _T_6464; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6466 = _T_6465 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6476 = _T_4726 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6477 = perr_ic_index_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6479 = _T_6477 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6480 = _T_6476 | _T_6479; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6481 = _T_6480 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6491 = _T_4727 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6492 = perr_ic_index_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6494 = _T_6492 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6495 = _T_6491 | _T_6494; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6496 = _T_6495 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6506 = _T_4728 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6507 = perr_ic_index_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6509 = _T_6507 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6510 = _T_6506 | _T_6509; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6511 = _T_6510 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6521 = _T_4729 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6522 = perr_ic_index_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6524 = _T_6522 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6525 = _T_6521 | _T_6524; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6526 = _T_6525 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6536 = _T_4730 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6537 = perr_ic_index_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6539 = _T_6537 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6540 = _T_6536 | _T_6539; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6541 = _T_6540 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6551 = _T_4731 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6552 = perr_ic_index_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6554 = _T_6552 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6555 = _T_6551 | _T_6554; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6556 = _T_6555 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6566 = _T_4732 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6567 = perr_ic_index_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6569 = _T_6567 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6570 = _T_6566 | _T_6569; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6571 = _T_6570 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6581 = _T_4733 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6582 = perr_ic_index_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_6584 = _T_6582 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6585 = _T_6581 | _T_6584; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6586 = _T_6585 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6596 = _T_4702 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6599 = _T_6117 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6600 = _T_6596 | _T_6599; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6601 = _T_6600 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6611 = _T_4703 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6614 = _T_6132 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6615 = _T_6611 | _T_6614; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6616 = _T_6615 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6626 = _T_4704 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6629 = _T_6147 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6630 = _T_6626 | _T_6629; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6631 = _T_6630 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6641 = _T_4705 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6644 = _T_6162 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6645 = _T_6641 | _T_6644; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6646 = _T_6645 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6656 = _T_4706 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6659 = _T_6177 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6660 = _T_6656 | _T_6659; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6661 = _T_6660 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6671 = _T_4707 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6674 = _T_6192 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6675 = _T_6671 | _T_6674; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6676 = _T_6675 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6686 = _T_4708 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6689 = _T_6207 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6690 = _T_6686 | _T_6689; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6691 = _T_6690 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6701 = _T_4709 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6704 = _T_6222 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6705 = _T_6701 | _T_6704; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6706 = _T_6705 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6716 = _T_4710 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6719 = _T_6237 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6720 = _T_6716 | _T_6719; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6721 = _T_6720 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6731 = _T_4711 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6734 = _T_6252 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6735 = _T_6731 | _T_6734; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6736 = _T_6735 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6746 = _T_4712 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6749 = _T_6267 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6750 = _T_6746 | _T_6749; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6751 = _T_6750 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6761 = _T_4713 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6764 = _T_6282 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6765 = _T_6761 | _T_6764; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6766 = _T_6765 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6776 = _T_4714 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6779 = _T_6297 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6780 = _T_6776 | _T_6779; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6781 = _T_6780 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6791 = _T_4715 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6794 = _T_6312 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6795 = _T_6791 | _T_6794; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6796 = _T_6795 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6806 = _T_4716 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6809 = _T_6327 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6810 = _T_6806 | _T_6809; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6811 = _T_6810 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6821 = _T_4717 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6824 = _T_6342 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6825 = _T_6821 | _T_6824; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6826 = _T_6825 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6836 = _T_4718 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6839 = _T_6357 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6840 = _T_6836 | _T_6839; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6841 = _T_6840 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6851 = _T_4719 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6854 = _T_6372 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6855 = _T_6851 | _T_6854; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6856 = _T_6855 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6866 = _T_4720 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6869 = _T_6387 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6870 = _T_6866 | _T_6869; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6871 = _T_6870 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6881 = _T_4721 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6884 = _T_6402 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6885 = _T_6881 | _T_6884; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6886 = _T_6885 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6896 = _T_4722 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6899 = _T_6417 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6900 = _T_6896 | _T_6899; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6901 = _T_6900 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6911 = _T_4723 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6914 = _T_6432 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6915 = _T_6911 | _T_6914; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6916 = _T_6915 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6926 = _T_4724 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6929 = _T_6447 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6930 = _T_6926 | _T_6929; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6931 = _T_6930 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6941 = _T_4725 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6944 = _T_6462 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6945 = _T_6941 | _T_6944; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6946 = _T_6945 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6956 = _T_4726 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6959 = _T_6477 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6960 = _T_6956 | _T_6959; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6961 = _T_6960 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6971 = _T_4727 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6974 = _T_6492 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6975 = _T_6971 | _T_6974; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6976 = _T_6975 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_6986 = _T_4728 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_6989 = _T_6507 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_6990 = _T_6986 | _T_6989; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_6991 = _T_6990 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7001 = _T_4729 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7004 = _T_6522 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7005 = _T_7001 | _T_7004; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7006 = _T_7005 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7016 = _T_4730 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7019 = _T_6537 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7020 = _T_7016 | _T_7019; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7021 = _T_7020 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7031 = _T_4731 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7034 = _T_6552 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7035 = _T_7031 | _T_7034; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7036 = _T_7035 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7046 = _T_4732 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7049 = _T_6567 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7050 = _T_7046 | _T_7049; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7051 = _T_7050 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7061 = _T_4733 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7064 = _T_6582 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7065 = _T_7061 | _T_7064; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7066 = _T_7065 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7076 = _T_4734 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7077 = perr_ic_index_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7079 = _T_7077 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7080 = _T_7076 | _T_7079; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7081 = _T_7080 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7091 = _T_4735 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7092 = perr_ic_index_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7094 = _T_7092 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7095 = _T_7091 | _T_7094; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7096 = _T_7095 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7106 = _T_4736 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7107 = perr_ic_index_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7109 = _T_7107 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7110 = _T_7106 | _T_7109; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7111 = _T_7110 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7121 = _T_4737 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7122 = perr_ic_index_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7124 = _T_7122 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7125 = _T_7121 | _T_7124; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7126 = _T_7125 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7136 = _T_4738 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7137 = perr_ic_index_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7139 = _T_7137 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7140 = _T_7136 | _T_7139; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7141 = _T_7140 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7151 = _T_4739 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7152 = perr_ic_index_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7154 = _T_7152 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7155 = _T_7151 | _T_7154; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7156 = _T_7155 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7166 = _T_4740 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7167 = perr_ic_index_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7169 = _T_7167 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7170 = _T_7166 | _T_7169; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7171 = _T_7170 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7181 = _T_4741 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7182 = perr_ic_index_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7184 = _T_7182 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7185 = _T_7181 | _T_7184; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7186 = _T_7185 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7196 = _T_4742 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7197 = perr_ic_index_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7199 = _T_7197 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7200 = _T_7196 | _T_7199; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7201 = _T_7200 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7211 = _T_4743 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7212 = perr_ic_index_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7214 = _T_7212 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7215 = _T_7211 | _T_7214; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7216 = _T_7215 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7226 = _T_4744 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7227 = perr_ic_index_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7229 = _T_7227 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7230 = _T_7226 | _T_7229; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7231 = _T_7230 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7241 = _T_4745 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7242 = perr_ic_index_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7244 = _T_7242 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7245 = _T_7241 | _T_7244; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7246 = _T_7245 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7256 = _T_4746 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7257 = perr_ic_index_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7259 = _T_7257 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7260 = _T_7256 | _T_7259; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7261 = _T_7260 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7271 = _T_4747 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7272 = perr_ic_index_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7274 = _T_7272 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7275 = _T_7271 | _T_7274; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7276 = _T_7275 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7286 = _T_4748 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7287 = perr_ic_index_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7289 = _T_7287 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7290 = _T_7286 | _T_7289; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7291 = _T_7290 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7301 = _T_4749 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7302 = perr_ic_index_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7304 = _T_7302 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7305 = _T_7301 | _T_7304; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7306 = _T_7305 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7316 = _T_4750 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7317 = perr_ic_index_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7319 = _T_7317 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7320 = _T_7316 | _T_7319; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7321 = _T_7320 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7331 = _T_4751 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7332 = perr_ic_index_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7334 = _T_7332 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7335 = _T_7331 | _T_7334; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7336 = _T_7335 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7346 = _T_4752 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7347 = perr_ic_index_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7349 = _T_7347 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7350 = _T_7346 | _T_7349; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7351 = _T_7350 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7361 = _T_4753 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7362 = perr_ic_index_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7364 = _T_7362 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7365 = _T_7361 | _T_7364; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7366 = _T_7365 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7376 = _T_4754 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7377 = perr_ic_index_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7379 = _T_7377 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7380 = _T_7376 | _T_7379; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7381 = _T_7380 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7391 = _T_4755 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7392 = perr_ic_index_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7394 = _T_7392 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7395 = _T_7391 | _T_7394; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7396 = _T_7395 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7406 = _T_4756 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7407 = perr_ic_index_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7409 = _T_7407 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7410 = _T_7406 | _T_7409; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7411 = _T_7410 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7421 = _T_4757 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7422 = perr_ic_index_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7424 = _T_7422 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7425 = _T_7421 | _T_7424; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7426 = _T_7425 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7436 = _T_4758 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7437 = perr_ic_index_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7439 = _T_7437 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7440 = _T_7436 | _T_7439; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7441 = _T_7440 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7451 = _T_4759 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7452 = perr_ic_index_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7454 = _T_7452 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7455 = _T_7451 | _T_7454; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7456 = _T_7455 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7466 = _T_4760 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7467 = perr_ic_index_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7469 = _T_7467 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7470 = _T_7466 | _T_7469; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7471 = _T_7470 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7481 = _T_4761 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7482 = perr_ic_index_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7484 = _T_7482 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7485 = _T_7481 | _T_7484; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7486 = _T_7485 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7496 = _T_4762 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7497 = perr_ic_index_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7499 = _T_7497 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7500 = _T_7496 | _T_7499; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7501 = _T_7500 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7511 = _T_4763 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7512 = perr_ic_index_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7514 = _T_7512 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7515 = _T_7511 | _T_7514; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7516 = _T_7515 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7526 = _T_4764 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7527 = perr_ic_index_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7529 = _T_7527 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7530 = _T_7526 | _T_7529; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7531 = _T_7530 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7541 = _T_4765 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7542 = perr_ic_index_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_7544 = _T_7542 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7545 = _T_7541 | _T_7544; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7546 = _T_7545 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7556 = _T_4734 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7559 = _T_7077 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7560 = _T_7556 | _T_7559; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7561 = _T_7560 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7571 = _T_4735 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7574 = _T_7092 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7575 = _T_7571 | _T_7574; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7576 = _T_7575 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7586 = _T_4736 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7589 = _T_7107 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7590 = _T_7586 | _T_7589; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7591 = _T_7590 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7601 = _T_4737 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7604 = _T_7122 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7605 = _T_7601 | _T_7604; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7606 = _T_7605 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7616 = _T_4738 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7619 = _T_7137 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7620 = _T_7616 | _T_7619; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7621 = _T_7620 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7631 = _T_4739 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7634 = _T_7152 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7635 = _T_7631 | _T_7634; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7636 = _T_7635 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7646 = _T_4740 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7649 = _T_7167 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7650 = _T_7646 | _T_7649; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7651 = _T_7650 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7661 = _T_4741 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7664 = _T_7182 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7665 = _T_7661 | _T_7664; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7666 = _T_7665 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7676 = _T_4742 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7679 = _T_7197 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7680 = _T_7676 | _T_7679; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7681 = _T_7680 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7691 = _T_4743 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7694 = _T_7212 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7695 = _T_7691 | _T_7694; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7696 = _T_7695 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7706 = _T_4744 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7709 = _T_7227 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7710 = _T_7706 | _T_7709; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7711 = _T_7710 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7721 = _T_4745 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7724 = _T_7242 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7725 = _T_7721 | _T_7724; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7726 = _T_7725 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7736 = _T_4746 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7739 = _T_7257 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7740 = _T_7736 | _T_7739; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7741 = _T_7740 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7751 = _T_4747 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7754 = _T_7272 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7755 = _T_7751 | _T_7754; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7756 = _T_7755 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7766 = _T_4748 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7769 = _T_7287 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7770 = _T_7766 | _T_7769; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7771 = _T_7770 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7781 = _T_4749 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7784 = _T_7302 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7785 = _T_7781 | _T_7784; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7786 = _T_7785 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7796 = _T_4750 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7799 = _T_7317 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7800 = _T_7796 | _T_7799; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7801 = _T_7800 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7811 = _T_4751 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7814 = _T_7332 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7815 = _T_7811 | _T_7814; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7816 = _T_7815 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7826 = _T_4752 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7829 = _T_7347 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7830 = _T_7826 | _T_7829; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7831 = _T_7830 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7841 = _T_4753 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7844 = _T_7362 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7845 = _T_7841 | _T_7844; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7846 = _T_7845 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7856 = _T_4754 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7859 = _T_7377 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7860 = _T_7856 | _T_7859; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7861 = _T_7860 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7871 = _T_4755 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7874 = _T_7392 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7875 = _T_7871 | _T_7874; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7876 = _T_7875 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7886 = _T_4756 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7889 = _T_7407 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7890 = _T_7886 | _T_7889; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7891 = _T_7890 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7901 = _T_4757 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7904 = _T_7422 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7905 = _T_7901 | _T_7904; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7906 = _T_7905 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7916 = _T_4758 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7919 = _T_7437 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7920 = _T_7916 | _T_7919; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7921 = _T_7920 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7931 = _T_4759 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7934 = _T_7452 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7935 = _T_7931 | _T_7934; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7936 = _T_7935 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7946 = _T_4760 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7949 = _T_7467 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7950 = _T_7946 | _T_7949; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7951 = _T_7950 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7961 = _T_4761 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7964 = _T_7482 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7965 = _T_7961 | _T_7964; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7966 = _T_7965 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7976 = _T_4762 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7979 = _T_7497 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7980 = _T_7976 | _T_7979; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7981 = _T_7980 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_7991 = _T_4763 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_7994 = _T_7512 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_7995 = _T_7991 | _T_7994; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_7996 = _T_7995 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8006 = _T_4764 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8009 = _T_7527 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8010 = _T_8006 | _T_8009; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8011 = _T_8010 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8021 = _T_4765 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8024 = _T_7542 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8025 = _T_8021 | _T_8024; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8026 = _T_8025 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8036 = _T_4766 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8037 = perr_ic_index_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8039 = _T_8037 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8040 = _T_8036 | _T_8039; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8041 = _T_8040 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8051 = _T_4767 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8052 = perr_ic_index_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8054 = _T_8052 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8055 = _T_8051 | _T_8054; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8056 = _T_8055 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8066 = _T_4768 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8067 = perr_ic_index_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8069 = _T_8067 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8070 = _T_8066 | _T_8069; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8071 = _T_8070 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8081 = _T_4769 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8082 = perr_ic_index_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8084 = _T_8082 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8085 = _T_8081 | _T_8084; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8086 = _T_8085 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8096 = _T_4770 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8097 = perr_ic_index_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8099 = _T_8097 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8100 = _T_8096 | _T_8099; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8101 = _T_8100 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8111 = _T_4771 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8112 = perr_ic_index_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8114 = _T_8112 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8115 = _T_8111 | _T_8114; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8116 = _T_8115 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8126 = _T_4772 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8127 = perr_ic_index_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8129 = _T_8127 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8130 = _T_8126 | _T_8129; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8131 = _T_8130 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8141 = _T_4773 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8142 = perr_ic_index_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8144 = _T_8142 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8145 = _T_8141 | _T_8144; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8146 = _T_8145 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8156 = _T_4774 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8157 = perr_ic_index_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8159 = _T_8157 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8160 = _T_8156 | _T_8159; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8161 = _T_8160 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8171 = _T_4775 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8172 = perr_ic_index_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8174 = _T_8172 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8175 = _T_8171 | _T_8174; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8176 = _T_8175 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8186 = _T_4776 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8187 = perr_ic_index_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8189 = _T_8187 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8190 = _T_8186 | _T_8189; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8191 = _T_8190 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8201 = _T_4777 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8202 = perr_ic_index_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8204 = _T_8202 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8205 = _T_8201 | _T_8204; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8206 = _T_8205 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8216 = _T_4778 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8217 = perr_ic_index_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8219 = _T_8217 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8220 = _T_8216 | _T_8219; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8221 = _T_8220 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8231 = _T_4779 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8232 = perr_ic_index_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8234 = _T_8232 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8235 = _T_8231 | _T_8234; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8236 = _T_8235 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8246 = _T_4780 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8247 = perr_ic_index_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8249 = _T_8247 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8250 = _T_8246 | _T_8249; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8251 = _T_8250 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8261 = _T_4781 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8262 = perr_ic_index_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8264 = _T_8262 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8265 = _T_8261 | _T_8264; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8266 = _T_8265 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8276 = _T_4782 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8277 = perr_ic_index_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8279 = _T_8277 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8280 = _T_8276 | _T_8279; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8281 = _T_8280 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8291 = _T_4783 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8292 = perr_ic_index_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8294 = _T_8292 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8295 = _T_8291 | _T_8294; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8296 = _T_8295 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8306 = _T_4784 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8307 = perr_ic_index_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8309 = _T_8307 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8310 = _T_8306 | _T_8309; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8311 = _T_8310 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8321 = _T_4785 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8322 = perr_ic_index_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8324 = _T_8322 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8325 = _T_8321 | _T_8324; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8326 = _T_8325 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8336 = _T_4786 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8337 = perr_ic_index_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8339 = _T_8337 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8340 = _T_8336 | _T_8339; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8341 = _T_8340 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8351 = _T_4787 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8352 = perr_ic_index_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8354 = _T_8352 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8355 = _T_8351 | _T_8354; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8356 = _T_8355 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8366 = _T_4788 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8367 = perr_ic_index_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8369 = _T_8367 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8370 = _T_8366 | _T_8369; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8371 = _T_8370 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8381 = _T_4789 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8382 = perr_ic_index_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8384 = _T_8382 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8385 = _T_8381 | _T_8384; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8386 = _T_8385 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8396 = _T_4790 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8397 = perr_ic_index_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8399 = _T_8397 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8400 = _T_8396 | _T_8399; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8401 = _T_8400 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8411 = _T_4791 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8412 = perr_ic_index_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8414 = _T_8412 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8415 = _T_8411 | _T_8414; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8416 = _T_8415 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8426 = _T_4792 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8427 = perr_ic_index_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8429 = _T_8427 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8430 = _T_8426 | _T_8429; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8431 = _T_8430 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8441 = _T_4793 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8442 = perr_ic_index_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8444 = _T_8442 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8445 = _T_8441 | _T_8444; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8446 = _T_8445 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8456 = _T_4794 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8457 = perr_ic_index_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8459 = _T_8457 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8460 = _T_8456 | _T_8459; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8461 = _T_8460 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8471 = _T_4795 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8472 = perr_ic_index_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8474 = _T_8472 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8475 = _T_8471 | _T_8474; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8476 = _T_8475 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8486 = _T_4796 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8487 = perr_ic_index_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8489 = _T_8487 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8490 = _T_8486 | _T_8489; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8491 = _T_8490 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8501 = _T_4797 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8502 = perr_ic_index_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 766:102]
  wire  _T_8504 = _T_8502 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8505 = _T_8501 | _T_8504; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8506 = _T_8505 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8516 = _T_4766 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8519 = _T_8037 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8520 = _T_8516 | _T_8519; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8521 = _T_8520 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8531 = _T_4767 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8534 = _T_8052 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8535 = _T_8531 | _T_8534; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8536 = _T_8535 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8546 = _T_4768 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8549 = _T_8067 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8550 = _T_8546 | _T_8549; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8551 = _T_8550 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8561 = _T_4769 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8564 = _T_8082 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8565 = _T_8561 | _T_8564; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8566 = _T_8565 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8576 = _T_4770 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8579 = _T_8097 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8580 = _T_8576 | _T_8579; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8581 = _T_8580 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8591 = _T_4771 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8594 = _T_8112 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8595 = _T_8591 | _T_8594; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8596 = _T_8595 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8606 = _T_4772 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8609 = _T_8127 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8610 = _T_8606 | _T_8609; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8611 = _T_8610 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8621 = _T_4773 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8624 = _T_8142 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8625 = _T_8621 | _T_8624; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8626 = _T_8625 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8636 = _T_4774 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8639 = _T_8157 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8640 = _T_8636 | _T_8639; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8641 = _T_8640 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8651 = _T_4775 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8654 = _T_8172 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8655 = _T_8651 | _T_8654; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8656 = _T_8655 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8666 = _T_4776 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8669 = _T_8187 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8670 = _T_8666 | _T_8669; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8671 = _T_8670 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8681 = _T_4777 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8684 = _T_8202 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8685 = _T_8681 | _T_8684; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8686 = _T_8685 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8696 = _T_4778 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8699 = _T_8217 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8700 = _T_8696 | _T_8699; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8701 = _T_8700 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8711 = _T_4779 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8714 = _T_8232 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8715 = _T_8711 | _T_8714; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8716 = _T_8715 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8726 = _T_4780 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8729 = _T_8247 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8730 = _T_8726 | _T_8729; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8731 = _T_8730 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8741 = _T_4781 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8744 = _T_8262 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8745 = _T_8741 | _T_8744; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8746 = _T_8745 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8756 = _T_4782 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8759 = _T_8277 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8760 = _T_8756 | _T_8759; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8761 = _T_8760 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8771 = _T_4783 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8774 = _T_8292 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8775 = _T_8771 | _T_8774; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8776 = _T_8775 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8786 = _T_4784 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8789 = _T_8307 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8790 = _T_8786 | _T_8789; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8791 = _T_8790 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8801 = _T_4785 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8804 = _T_8322 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8805 = _T_8801 | _T_8804; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8806 = _T_8805 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8816 = _T_4786 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8819 = _T_8337 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8820 = _T_8816 | _T_8819; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8821 = _T_8820 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8831 = _T_4787 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8834 = _T_8352 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8835 = _T_8831 | _T_8834; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8836 = _T_8835 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8846 = _T_4788 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8849 = _T_8367 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8850 = _T_8846 | _T_8849; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8851 = _T_8850 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8861 = _T_4789 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8864 = _T_8382 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8865 = _T_8861 | _T_8864; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8866 = _T_8865 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8876 = _T_4790 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8879 = _T_8397 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8880 = _T_8876 | _T_8879; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8881 = _T_8880 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8891 = _T_4791 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8894 = _T_8412 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8895 = _T_8891 | _T_8894; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8896 = _T_8895 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8906 = _T_4792 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8909 = _T_8427 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8910 = _T_8906 | _T_8909; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8911 = _T_8910 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8921 = _T_4793 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8924 = _T_8442 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8925 = _T_8921 | _T_8924; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8926 = _T_8925 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8936 = _T_4794 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8939 = _T_8457 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8940 = _T_8936 | _T_8939; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8941 = _T_8940 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8951 = _T_4795 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8954 = _T_8472 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8955 = _T_8951 | _T_8954; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8956 = _T_8955 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8966 = _T_4796 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8969 = _T_8487 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8970 = _T_8966 | _T_8969; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8971 = _T_8970 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_8981 = _T_4797 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 766:59]
  wire  _T_8984 = _T_8502 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 766:124]
  wire  _T_8985 = _T_8981 | _T_8984; // @[el2_ifu_mem_ctl.scala 766:81]
  wire  _T_8986 = _T_8985 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 766:147]
  wire  _T_9788 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 821:63]
  wire  _T_9789 = _T_9788 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 821:85]
  wire [1:0] _T_9791 = _T_9789 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_9798; // @[el2_ifu_mem_ctl.scala 826:57]
  reg  _T_9799; // @[el2_ifu_mem_ctl.scala 827:56]
  reg  _T_9800; // @[el2_ifu_mem_ctl.scala 828:59]
  wire  _T_9801 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 829:80]
  wire  _T_9802 = ifu_bus_arvalid_ff & _T_9801; // @[el2_ifu_mem_ctl.scala 829:78]
  reg  _T_9804; // @[el2_ifu_mem_ctl.scala 829:58]
  reg  _T_9805; // @[el2_ifu_mem_ctl.scala 830:58]
  wire  _T_9808 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 837:71]
  wire  _T_9810 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 837:124]
  wire  _T_9812 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 838:50]
  wire  _T_9814 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 838:103]
  wire [3:0] _T_9817 = {_T_9808,_T_9810,_T_9812,_T_9814}; // @[Cat.scala 29:58]
  reg  _T_9826; // @[Reg.scala 27:20]
  wire [31:0] _T_9836 = {io_ifc_fetch_addr_bf,1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_9837 = _T_9836 | 32'h7fffffff; // @[el2_ifu_mem_ctl.scala 846:65]
  wire  _T_9839 = _T_9837 == 32'h7fffffff; // @[el2_ifu_mem_ctl.scala 846:96]
  wire [31:0] _T_9843 = _T_9836 | 32'h3fffffff; // @[el2_ifu_mem_ctl.scala 847:65]
  wire  _T_9845 = _T_9843 == 32'hffffffff; // @[el2_ifu_mem_ctl.scala 847:96]
  wire  _T_9847 = _T_9839 | _T_9845; // @[el2_ifu_mem_ctl.scala 846:162]
  wire [31:0] _T_9849 = _T_9836 | 32'h1fffffff; // @[el2_ifu_mem_ctl.scala 848:65]
  wire  _T_9851 = _T_9849 == 32'hbfffffff; // @[el2_ifu_mem_ctl.scala 848:96]
  wire  _T_9853 = _T_9847 | _T_9851; // @[el2_ifu_mem_ctl.scala 847:162]
  wire [31:0] _T_9855 = _T_9836 | 32'hfffffff; // @[el2_ifu_mem_ctl.scala 849:65]
  wire  _T_9857 = _T_9855 == 32'h8fffffff; // @[el2_ifu_mem_ctl.scala 849:96]
  wire  ifc_region_acc_okay = _T_9853 | _T_9857; // @[el2_ifu_mem_ctl.scala 848:162]
  wire  _T_9884 = ~ifc_region_acc_okay; // @[el2_ifu_mem_ctl.scala 854:65]
  wire  _T_9885 = _T_3938 & _T_9884; // @[el2_ifu_mem_ctl.scala 854:63]
  wire  ifc_region_acc_fault_memory_bf = _T_9885 & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 854:86]
  rvclkhdr rvclkhdr ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  rvclkhdr rvclkhdr_26 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_26_io_l1clk),
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en),
    .io_scan_mode(rvclkhdr_26_io_scan_mode)
  );
  rvclkhdr rvclkhdr_27 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_27_io_l1clk),
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en),
    .io_scan_mode(rvclkhdr_27_io_scan_mode)
  );
  rvclkhdr rvclkhdr_28 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_28_io_l1clk),
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en),
    .io_scan_mode(rvclkhdr_28_io_scan_mode)
  );
  rvclkhdr rvclkhdr_29 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_29_io_l1clk),
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en),
    .io_scan_mode(rvclkhdr_29_io_scan_mode)
  );
  rvclkhdr rvclkhdr_30 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_30_io_l1clk),
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en),
    .io_scan_mode(rvclkhdr_30_io_scan_mode)
  );
  rvclkhdr rvclkhdr_31 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_31_io_l1clk),
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en),
    .io_scan_mode(rvclkhdr_31_io_scan_mode)
  );
  rvclkhdr rvclkhdr_32 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_32_io_l1clk),
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en),
    .io_scan_mode(rvclkhdr_32_io_scan_mode)
  );
  rvclkhdr rvclkhdr_33 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_33_io_l1clk),
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en),
    .io_scan_mode(rvclkhdr_33_io_scan_mode)
  );
  rvclkhdr rvclkhdr_34 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_34_io_l1clk),
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en),
    .io_scan_mode(rvclkhdr_34_io_scan_mode)
  );
  rvclkhdr rvclkhdr_35 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_35_io_l1clk),
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en),
    .io_scan_mode(rvclkhdr_35_io_scan_mode)
  );
  rvclkhdr rvclkhdr_36 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_36_io_l1clk),
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en),
    .io_scan_mode(rvclkhdr_36_io_scan_mode)
  );
  rvclkhdr rvclkhdr_37 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_37_io_l1clk),
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en),
    .io_scan_mode(rvclkhdr_37_io_scan_mode)
  );
  rvclkhdr rvclkhdr_38 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_38_io_l1clk),
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en),
    .io_scan_mode(rvclkhdr_38_io_scan_mode)
  );
  rvclkhdr rvclkhdr_39 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_39_io_l1clk),
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en),
    .io_scan_mode(rvclkhdr_39_io_scan_mode)
  );
  rvclkhdr rvclkhdr_40 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_40_io_l1clk),
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en),
    .io_scan_mode(rvclkhdr_40_io_scan_mode)
  );
  rvclkhdr rvclkhdr_41 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_41_io_l1clk),
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en),
    .io_scan_mode(rvclkhdr_41_io_scan_mode)
  );
  rvclkhdr rvclkhdr_42 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_42_io_l1clk),
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en),
    .io_scan_mode(rvclkhdr_42_io_scan_mode)
  );
  rvclkhdr rvclkhdr_43 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_43_io_l1clk),
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en),
    .io_scan_mode(rvclkhdr_43_io_scan_mode)
  );
  rvclkhdr rvclkhdr_44 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_44_io_l1clk),
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en),
    .io_scan_mode(rvclkhdr_44_io_scan_mode)
  );
  rvclkhdr rvclkhdr_45 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_45_io_l1clk),
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en),
    .io_scan_mode(rvclkhdr_45_io_scan_mode)
  );
  rvclkhdr rvclkhdr_46 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_46_io_l1clk),
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en),
    .io_scan_mode(rvclkhdr_46_io_scan_mode)
  );
  rvclkhdr rvclkhdr_47 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_47_io_l1clk),
    .io_clk(rvclkhdr_47_io_clk),
    .io_en(rvclkhdr_47_io_en),
    .io_scan_mode(rvclkhdr_47_io_scan_mode)
  );
  rvclkhdr rvclkhdr_48 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_48_io_l1clk),
    .io_clk(rvclkhdr_48_io_clk),
    .io_en(rvclkhdr_48_io_en),
    .io_scan_mode(rvclkhdr_48_io_scan_mode)
  );
  rvclkhdr rvclkhdr_49 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_49_io_l1clk),
    .io_clk(rvclkhdr_49_io_clk),
    .io_en(rvclkhdr_49_io_en),
    .io_scan_mode(rvclkhdr_49_io_scan_mode)
  );
  rvclkhdr rvclkhdr_50 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_50_io_l1clk),
    .io_clk(rvclkhdr_50_io_clk),
    .io_en(rvclkhdr_50_io_en),
    .io_scan_mode(rvclkhdr_50_io_scan_mode)
  );
  rvclkhdr rvclkhdr_51 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_51_io_l1clk),
    .io_clk(rvclkhdr_51_io_clk),
    .io_en(rvclkhdr_51_io_en),
    .io_scan_mode(rvclkhdr_51_io_scan_mode)
  );
  rvclkhdr rvclkhdr_52 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_52_io_l1clk),
    .io_clk(rvclkhdr_52_io_clk),
    .io_en(rvclkhdr_52_io_en),
    .io_scan_mode(rvclkhdr_52_io_scan_mode)
  );
  rvclkhdr rvclkhdr_53 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_53_io_l1clk),
    .io_clk(rvclkhdr_53_io_clk),
    .io_en(rvclkhdr_53_io_en),
    .io_scan_mode(rvclkhdr_53_io_scan_mode)
  );
  rvclkhdr rvclkhdr_54 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_54_io_l1clk),
    .io_clk(rvclkhdr_54_io_clk),
    .io_en(rvclkhdr_54_io_en),
    .io_scan_mode(rvclkhdr_54_io_scan_mode)
  );
  rvclkhdr rvclkhdr_55 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_55_io_l1clk),
    .io_clk(rvclkhdr_55_io_clk),
    .io_en(rvclkhdr_55_io_en),
    .io_scan_mode(rvclkhdr_55_io_scan_mode)
  );
  rvclkhdr rvclkhdr_56 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_56_io_l1clk),
    .io_clk(rvclkhdr_56_io_clk),
    .io_en(rvclkhdr_56_io_en),
    .io_scan_mode(rvclkhdr_56_io_scan_mode)
  );
  rvclkhdr rvclkhdr_57 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_57_io_l1clk),
    .io_clk(rvclkhdr_57_io_clk),
    .io_en(rvclkhdr_57_io_en),
    .io_scan_mode(rvclkhdr_57_io_scan_mode)
  );
  rvclkhdr rvclkhdr_58 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_58_io_l1clk),
    .io_clk(rvclkhdr_58_io_clk),
    .io_en(rvclkhdr_58_io_en),
    .io_scan_mode(rvclkhdr_58_io_scan_mode)
  );
  rvclkhdr rvclkhdr_59 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_59_io_l1clk),
    .io_clk(rvclkhdr_59_io_clk),
    .io_en(rvclkhdr_59_io_en),
    .io_scan_mode(rvclkhdr_59_io_scan_mode)
  );
  rvclkhdr rvclkhdr_60 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_60_io_l1clk),
    .io_clk(rvclkhdr_60_io_clk),
    .io_en(rvclkhdr_60_io_en),
    .io_scan_mode(rvclkhdr_60_io_scan_mode)
  );
  rvclkhdr rvclkhdr_61 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_61_io_l1clk),
    .io_clk(rvclkhdr_61_io_clk),
    .io_en(rvclkhdr_61_io_en),
    .io_scan_mode(rvclkhdr_61_io_scan_mode)
  );
  rvclkhdr rvclkhdr_62 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_62_io_l1clk),
    .io_clk(rvclkhdr_62_io_clk),
    .io_en(rvclkhdr_62_io_en),
    .io_scan_mode(rvclkhdr_62_io_scan_mode)
  );
  rvclkhdr rvclkhdr_63 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_63_io_l1clk),
    .io_clk(rvclkhdr_63_io_clk),
    .io_en(rvclkhdr_63_io_en),
    .io_scan_mode(rvclkhdr_63_io_scan_mode)
  );
  rvclkhdr rvclkhdr_64 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_64_io_l1clk),
    .io_clk(rvclkhdr_64_io_clk),
    .io_en(rvclkhdr_64_io_en),
    .io_scan_mode(rvclkhdr_64_io_scan_mode)
  );
  rvclkhdr rvclkhdr_65 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_65_io_l1clk),
    .io_clk(rvclkhdr_65_io_clk),
    .io_en(rvclkhdr_65_io_en),
    .io_scan_mode(rvclkhdr_65_io_scan_mode)
  );
  rvclkhdr rvclkhdr_66 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_66_io_l1clk),
    .io_clk(rvclkhdr_66_io_clk),
    .io_en(rvclkhdr_66_io_en),
    .io_scan_mode(rvclkhdr_66_io_scan_mode)
  );
  rvclkhdr rvclkhdr_67 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_67_io_l1clk),
    .io_clk(rvclkhdr_67_io_clk),
    .io_en(rvclkhdr_67_io_en),
    .io_scan_mode(rvclkhdr_67_io_scan_mode)
  );
  rvclkhdr rvclkhdr_68 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_68_io_l1clk),
    .io_clk(rvclkhdr_68_io_clk),
    .io_en(rvclkhdr_68_io_en),
    .io_scan_mode(rvclkhdr_68_io_scan_mode)
  );
  rvclkhdr rvclkhdr_69 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_69_io_l1clk),
    .io_clk(rvclkhdr_69_io_clk),
    .io_en(rvclkhdr_69_io_en),
    .io_scan_mode(rvclkhdr_69_io_scan_mode)
  );
  rvclkhdr rvclkhdr_70 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_70_io_l1clk),
    .io_clk(rvclkhdr_70_io_clk),
    .io_en(rvclkhdr_70_io_en),
    .io_scan_mode(rvclkhdr_70_io_scan_mode)
  );
  rvclkhdr rvclkhdr_71 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_71_io_l1clk),
    .io_clk(rvclkhdr_71_io_clk),
    .io_en(rvclkhdr_71_io_en),
    .io_scan_mode(rvclkhdr_71_io_scan_mode)
  );
  rvclkhdr rvclkhdr_72 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_72_io_l1clk),
    .io_clk(rvclkhdr_72_io_clk),
    .io_en(rvclkhdr_72_io_en),
    .io_scan_mode(rvclkhdr_72_io_scan_mode)
  );
  rvclkhdr rvclkhdr_73 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_73_io_l1clk),
    .io_clk(rvclkhdr_73_io_clk),
    .io_en(rvclkhdr_73_io_en),
    .io_scan_mode(rvclkhdr_73_io_scan_mode)
  );
  rvclkhdr rvclkhdr_74 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_74_io_l1clk),
    .io_clk(rvclkhdr_74_io_clk),
    .io_en(rvclkhdr_74_io_en),
    .io_scan_mode(rvclkhdr_74_io_scan_mode)
  );
  rvclkhdr rvclkhdr_75 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_75_io_l1clk),
    .io_clk(rvclkhdr_75_io_clk),
    .io_en(rvclkhdr_75_io_en),
    .io_scan_mode(rvclkhdr_75_io_scan_mode)
  );
  rvclkhdr rvclkhdr_76 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_76_io_l1clk),
    .io_clk(rvclkhdr_76_io_clk),
    .io_en(rvclkhdr_76_io_en),
    .io_scan_mode(rvclkhdr_76_io_scan_mode)
  );
  rvclkhdr rvclkhdr_77 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_77_io_l1clk),
    .io_clk(rvclkhdr_77_io_clk),
    .io_en(rvclkhdr_77_io_en),
    .io_scan_mode(rvclkhdr_77_io_scan_mode)
  );
  rvclkhdr rvclkhdr_78 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_78_io_l1clk),
    .io_clk(rvclkhdr_78_io_clk),
    .io_en(rvclkhdr_78_io_en),
    .io_scan_mode(rvclkhdr_78_io_scan_mode)
  );
  rvclkhdr rvclkhdr_79 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_79_io_l1clk),
    .io_clk(rvclkhdr_79_io_clk),
    .io_en(rvclkhdr_79_io_en),
    .io_scan_mode(rvclkhdr_79_io_scan_mode)
  );
  rvclkhdr rvclkhdr_80 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_80_io_l1clk),
    .io_clk(rvclkhdr_80_io_clk),
    .io_en(rvclkhdr_80_io_en),
    .io_scan_mode(rvclkhdr_80_io_scan_mode)
  );
  rvclkhdr rvclkhdr_81 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_81_io_l1clk),
    .io_clk(rvclkhdr_81_io_clk),
    .io_en(rvclkhdr_81_io_en),
    .io_scan_mode(rvclkhdr_81_io_scan_mode)
  );
  rvclkhdr rvclkhdr_82 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_82_io_l1clk),
    .io_clk(rvclkhdr_82_io_clk),
    .io_en(rvclkhdr_82_io_en),
    .io_scan_mode(rvclkhdr_82_io_scan_mode)
  );
  rvclkhdr rvclkhdr_83 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_83_io_l1clk),
    .io_clk(rvclkhdr_83_io_clk),
    .io_en(rvclkhdr_83_io_en),
    .io_scan_mode(rvclkhdr_83_io_scan_mode)
  );
  rvclkhdr rvclkhdr_84 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_84_io_l1clk),
    .io_clk(rvclkhdr_84_io_clk),
    .io_en(rvclkhdr_84_io_en),
    .io_scan_mode(rvclkhdr_84_io_scan_mode)
  );
  rvclkhdr rvclkhdr_85 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_85_io_l1clk),
    .io_clk(rvclkhdr_85_io_clk),
    .io_en(rvclkhdr_85_io_en),
    .io_scan_mode(rvclkhdr_85_io_scan_mode)
  );
  rvclkhdr rvclkhdr_86 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_86_io_l1clk),
    .io_clk(rvclkhdr_86_io_clk),
    .io_en(rvclkhdr_86_io_en),
    .io_scan_mode(rvclkhdr_86_io_scan_mode)
  );
  rvclkhdr rvclkhdr_87 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_87_io_l1clk),
    .io_clk(rvclkhdr_87_io_clk),
    .io_en(rvclkhdr_87_io_en),
    .io_scan_mode(rvclkhdr_87_io_scan_mode)
  );
  rvclkhdr rvclkhdr_88 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_88_io_l1clk),
    .io_clk(rvclkhdr_88_io_clk),
    .io_en(rvclkhdr_88_io_en),
    .io_scan_mode(rvclkhdr_88_io_scan_mode)
  );
  rvclkhdr rvclkhdr_89 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_89_io_l1clk),
    .io_clk(rvclkhdr_89_io_clk),
    .io_en(rvclkhdr_89_io_en),
    .io_scan_mode(rvclkhdr_89_io_scan_mode)
  );
  rvclkhdr rvclkhdr_90 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_90_io_l1clk),
    .io_clk(rvclkhdr_90_io_clk),
    .io_en(rvclkhdr_90_io_en),
    .io_scan_mode(rvclkhdr_90_io_scan_mode)
  );
  rvclkhdr rvclkhdr_91 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_91_io_l1clk),
    .io_clk(rvclkhdr_91_io_clk),
    .io_en(rvclkhdr_91_io_en),
    .io_scan_mode(rvclkhdr_91_io_scan_mode)
  );
  rvclkhdr rvclkhdr_92 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_92_io_l1clk),
    .io_clk(rvclkhdr_92_io_clk),
    .io_en(rvclkhdr_92_io_en),
    .io_scan_mode(rvclkhdr_92_io_scan_mode)
  );
  rvclkhdr rvclkhdr_93 ( // @[el2_lib.scala 483:22]
    .io_l1clk(rvclkhdr_93_io_l1clk),
    .io_clk(rvclkhdr_93_io_clk),
    .io_en(rvclkhdr_93_io_en),
    .io_scan_mode(rvclkhdr_93_io_scan_mode)
  );
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 330:26]
  assign io_ifu_ic_mb_empty = _T_328 | _T_231; // @[el2_ifu_mem_ctl.scala 329:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 193:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3987; // @[el2_ifu_mem_ctl.scala 709:21]
  assign io_ifu_pmu_ic_miss = _T_9798; // @[el2_ifu_mem_ctl.scala 826:22]
  assign io_ifu_pmu_ic_hit = _T_9799; // @[el2_ifu_mem_ctl.scala 827:21]
  assign io_ifu_pmu_bus_error = _T_9800; // @[el2_ifu_mem_ctl.scala 828:24]
  assign io_ifu_pmu_bus_busy = _T_9804; // @[el2_ifu_mem_ctl.scala 829:23]
  assign io_ifu_pmu_bus_trxn = _T_9805; // @[el2_ifu_mem_ctl.scala 830:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 144:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 143:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 138:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 142:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 140:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 151:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 153:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 148:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 146:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 139:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 137:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 135:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 136:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 145:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 154:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 149:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 570:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2607; // @[el2_ifu_mem_ctl.scala 571:19]
  assign io_ifu_axi_araddr = _T_2609 & _T_2611; // @[el2_ifu_mem_ctl.scala 572:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 575:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 150:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 573:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 576:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 141:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 574:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 152:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 147:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 577:21]
  assign io_iccm_dma_ecc_error = iccm_dma_ecc_error; // @[el2_ifu_mem_ctl.scala 668:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 666:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 670:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 661:20]
  assign io_iccm_ready = _T_2705 & _T_2699; // @[el2_ifu_mem_ctl.scala 640:17]
  assign io_ic_rw_addr = _T_340 | _T_341; // @[el2_ifu_mem_ctl.scala 339:17]
  assign io_ic_wr_en = bus_ic_wr_en & _T_3973; // @[el2_ifu_mem_ctl.scala 708:15]
  assign io_ic_rd_en = _T_3965 | _T_3970; // @[el2_ifu_mem_ctl.scala 699:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 346:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 346:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 347:23]
  assign io_ifu_ic_debug_rd_data = _T_1211; // @[el2_ifu_mem_ctl.scala 355:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 833:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 835:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 836:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 834:25]
  assign io_ic_debug_way = _T_9817[1:0]; // @[el2_ifu_mem_ctl.scala 837:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_9791; // @[el2_ifu_mem_ctl.scala 821:19]
  assign io_iccm_rw_addr = _T_3109 ? io_dma_mem_addr[15:1] : _T_3116; // @[el2_ifu_mem_ctl.scala 672:19]
  assign io_iccm_wren = _T_2709 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 642:16]
  assign io_iccm_rden = _T_2713 | _T_2714; // @[el2_ifu_mem_ctl.scala 643:16]
  assign io_iccm_wr_data = _T_3091 ? _T_3092 : _T_3099; // @[el2_ifu_mem_ctl.scala 649:19]
  assign io_iccm_wr_size = _T_2719 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 645:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 290:15]
  assign io_ic_access_fault_f = _T_2491 & _T_319; // @[el2_ifu_mem_ctl.scala 393:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1277; // @[el2_ifu_mem_ctl.scala 394:29]
  assign io_iccm_rd_ecc_single_err = _T_3910 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 685:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 686:29]
  assign io_ic_error_start = _T_1199 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 349:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 192:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 191:24]
  assign io_ic_fetch_val_f = {_T_1285,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 397:21]
  assign io_ic_data_f = ic_final_data[31:0]; // @[el2_ifu_mem_ctl.scala 390:16]
  assign io_ic_premux_data = ic_premux_data_temp[63:0]; // @[el2_ifu_mem_ctl.scala 387:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 388:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_9826; // @[el2_ifu_mem_ctl.scala 844:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2496; // @[el2_ifu_mem_ctl.scala 487:27]
  assign io_iccm_correction_state = _T_2525 ? 1'h0 : _GEN_42; // @[el2_ifu_mem_ctl.scala 522:28 el2_ifu_mem_ctl.scala 535:32 el2_ifu_mem_ctl.scala 542:32 el2_ifu_mem_ctl.scala 549:32]
  assign rvclkhdr_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_io_en = ic_debug_rd_en_ff; // @[el2_lib.scala 485:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_1_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_1_io_en = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_lib.scala 485:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_2_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_2_io_en = _T_2 | scnd_miss_req; // @[el2_lib.scala 485:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_3_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_3_io_en = _T_309 | io_dec_tlu_force_halt; // @[el2_lib.scala 485:16]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_4_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_4_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_5_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_5_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_6_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_6_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_7_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_7_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_8_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_8_io_en = bus_ifu_wr_en & _T_1292; // @[el2_lib.scala 485:16]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_9_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_9_io_en = bus_ifu_wr_en & _T_1293; // @[el2_lib.scala 485:16]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_10_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_10_io_en = bus_ifu_wr_en & _T_1294; // @[el2_lib.scala 485:16]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_11_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_11_io_en = bus_ifu_wr_en & _T_1295; // @[el2_lib.scala 485:16]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_12_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_12_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_13_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_13_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_14_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_14_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_15_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_15_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_16_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_16_io_en = bus_ifu_wr_en & _T_1292; // @[el2_lib.scala 485:16]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_17_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_17_io_en = bus_ifu_wr_en & _T_1293; // @[el2_lib.scala 485:16]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_18_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_18_io_en = bus_ifu_wr_en & _T_1294; // @[el2_lib.scala 485:16]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_19_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_19_io_en = bus_ifu_wr_en & _T_1295; // @[el2_lib.scala 485:16]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_20_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_20_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_21_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_21_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_22_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_22_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_23_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_23_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_24_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_24_io_en = bus_ifu_wr_en & _T_1292; // @[el2_lib.scala 485:16]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_25_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_25_io_en = bus_ifu_wr_en & _T_1293; // @[el2_lib.scala 485:16]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_26_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_26_io_en = bus_ifu_wr_en & _T_1294; // @[el2_lib.scala 485:16]
  assign rvclkhdr_26_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_27_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_27_io_en = bus_ifu_wr_en & _T_1295; // @[el2_lib.scala 485:16]
  assign rvclkhdr_27_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_28_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_28_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_28_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_29_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_29_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_29_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_30_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_30_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_30_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_31_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_31_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_31_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_32_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_32_io_en = bus_ifu_wr_en & _T_1292; // @[el2_lib.scala 485:16]
  assign rvclkhdr_32_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_33_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_33_io_en = bus_ifu_wr_en & _T_1293; // @[el2_lib.scala 485:16]
  assign rvclkhdr_33_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_34_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_34_io_en = bus_ifu_wr_en & _T_1294; // @[el2_lib.scala 485:16]
  assign rvclkhdr_34_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_35_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_35_io_en = bus_ifu_wr_en & _T_1295; // @[el2_lib.scala 485:16]
  assign rvclkhdr_35_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_36_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_36_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_36_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_37_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_37_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_37_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_38_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_38_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_38_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_39_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_39_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_39_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_40_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_40_io_en = bus_ifu_wr_en & _T_1292; // @[el2_lib.scala 485:16]
  assign rvclkhdr_40_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_41_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_41_io_en = bus_ifu_wr_en & _T_1293; // @[el2_lib.scala 485:16]
  assign rvclkhdr_41_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_42_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_42_io_en = bus_ifu_wr_en & _T_1294; // @[el2_lib.scala 485:16]
  assign rvclkhdr_42_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_43_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_43_io_en = bus_ifu_wr_en & _T_1295; // @[el2_lib.scala 485:16]
  assign rvclkhdr_43_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_44_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_44_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_44_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_45_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_45_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_45_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_46_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_46_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_46_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_47_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_47_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_47_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_48_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_48_io_en = bus_ifu_wr_en & _T_1292; // @[el2_lib.scala 485:16]
  assign rvclkhdr_48_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_49_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_49_io_en = bus_ifu_wr_en & _T_1293; // @[el2_lib.scala 485:16]
  assign rvclkhdr_49_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_50_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_50_io_en = bus_ifu_wr_en & _T_1294; // @[el2_lib.scala 485:16]
  assign rvclkhdr_50_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_51_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_51_io_en = bus_ifu_wr_en & _T_1295; // @[el2_lib.scala 485:16]
  assign rvclkhdr_51_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_52_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_52_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_52_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_53_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_53_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_53_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_54_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_54_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_54_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_55_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_55_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_55_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_56_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_56_io_en = bus_ifu_wr_en & _T_1292; // @[el2_lib.scala 485:16]
  assign rvclkhdr_56_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_57_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_57_io_en = bus_ifu_wr_en & _T_1293; // @[el2_lib.scala 485:16]
  assign rvclkhdr_57_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_58_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_58_io_en = bus_ifu_wr_en & _T_1294; // @[el2_lib.scala 485:16]
  assign rvclkhdr_58_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_59_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_59_io_en = bus_ifu_wr_en & _T_1295; // @[el2_lib.scala 485:16]
  assign rvclkhdr_59_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_60_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_60_io_en = bus_ifu_wr_en & _T_1288; // @[el2_lib.scala 485:16]
  assign rvclkhdr_60_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_61_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_61_io_en = bus_ifu_wr_en & _T_1289; // @[el2_lib.scala 485:16]
  assign rvclkhdr_61_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_62_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_62_io_en = bus_ifu_wr_en & _T_1290; // @[el2_lib.scala 485:16]
  assign rvclkhdr_62_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_63_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_63_io_en = bus_ifu_wr_en & _T_1291; // @[el2_lib.scala 485:16]
  assign rvclkhdr_63_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_64_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_64_io_en = bus_ifu_wr_en & _T_1292; // @[el2_lib.scala 485:16]
  assign rvclkhdr_64_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_65_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_65_io_en = bus_ifu_wr_en & _T_1293; // @[el2_lib.scala 485:16]
  assign rvclkhdr_65_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_66_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_66_io_en = bus_ifu_wr_en & _T_1294; // @[el2_lib.scala 485:16]
  assign rvclkhdr_66_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_67_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_67_io_en = bus_ifu_wr_en & _T_1295; // @[el2_lib.scala 485:16]
  assign rvclkhdr_67_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_68_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_68_io_en = io_ifu_bus_clk_en; // @[el2_lib.scala 485:16]
  assign rvclkhdr_68_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_69_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_69_io_en = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_lib.scala 485:16]
  assign rvclkhdr_69_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_70_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_70_io_en = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_lib.scala 485:16]
  assign rvclkhdr_70_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_71_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_71_io_en = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_lib.scala 485:16]
  assign rvclkhdr_71_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_72_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_72_io_en = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_lib.scala 485:16]
  assign rvclkhdr_72_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_73_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_73_io_en = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_lib.scala 485:16]
  assign rvclkhdr_73_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_74_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_74_io_en = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_lib.scala 485:16]
  assign rvclkhdr_74_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_75_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_75_io_en = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_lib.scala 485:16]
  assign rvclkhdr_75_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_76_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_76_io_en = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_lib.scala 485:16]
  assign rvclkhdr_76_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_77_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_77_io_en = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_lib.scala 485:16]
  assign rvclkhdr_77_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_78_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_78_io_en = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_lib.scala 485:16]
  assign rvclkhdr_78_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_79_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_79_io_en = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_lib.scala 485:16]
  assign rvclkhdr_79_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_80_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_80_io_en = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_lib.scala 485:16]
  assign rvclkhdr_80_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_81_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_81_io_en = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_lib.scala 485:16]
  assign rvclkhdr_81_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_82_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_82_io_en = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_lib.scala 485:16]
  assign rvclkhdr_82_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_83_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_83_io_en = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_lib.scala 485:16]
  assign rvclkhdr_83_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_84_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_84_io_en = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_lib.scala 485:16]
  assign rvclkhdr_84_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_85_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_85_io_en = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_lib.scala 485:16]
  assign rvclkhdr_85_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_86_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_86_io_en = tag_valid_clken_0[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_86_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_87_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_87_io_en = tag_valid_clken_0[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_87_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_88_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_88_io_en = tag_valid_clken_1[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_88_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_89_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_89_io_en = tag_valid_clken_1[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_89_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_90_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_90_io_en = tag_valid_clken_2[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_90_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_91_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_91_io_en = tag_valid_clken_2[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_91_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_92_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_92_io_en = tag_valid_clken_3[0]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_92_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
  assign rvclkhdr_93_io_clk = clock; // @[el2_lib.scala 484:17]
  assign rvclkhdr_93_io_en = tag_valid_clken_3[1]; // @[el2_lib.scala 485:16]
  assign rvclkhdr_93_io_scan_mode = io_scan_mode; // @[el2_lib.scala 486:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ifu_ic_rw_int_addr_ff = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  way_status_out_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_status_out_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_status_out_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_status_out_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_status_out_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_status_out_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_status_out_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_status_out_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_status_out_8 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_status_out_9 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_status_out_10 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_status_out_11 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_status_out_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_status_out_13 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_status_out_14 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_status_out_15 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_status_out_16 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_status_out_17 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_status_out_18 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_status_out_19 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_status_out_20 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_status_out_21 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_status_out_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_status_out_23 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_status_out_24 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_status_out_25 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_status_out_26 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_status_out_27 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_status_out_28 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_status_out_29 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_status_out_30 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_status_out_31 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_status_out_32 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_status_out_33 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_status_out_34 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_status_out_35 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_status_out_36 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_status_out_37 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_status_out_38 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_status_out_39 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_status_out_40 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_status_out_41 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way_status_out_42 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way_status_out_43 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way_status_out_44 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way_status_out_45 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way_status_out_46 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way_status_out_47 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way_status_out_48 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way_status_out_49 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way_status_out_50 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way_status_out_51 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way_status_out_52 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way_status_out_53 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way_status_out_54 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way_status_out_55 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way_status_out_56 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way_status_out_57 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way_status_out_58 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way_status_out_59 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way_status_out_60 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way_status_out_61 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way_status_out_62 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way_status_out_63 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way_status_out_64 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way_status_out_65 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way_status_out_66 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way_status_out_67 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way_status_out_68 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way_status_out_69 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way_status_out_70 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way_status_out_71 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way_status_out_72 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way_status_out_73 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way_status_out_74 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way_status_out_75 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way_status_out_76 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way_status_out_77 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way_status_out_78 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way_status_out_79 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way_status_out_80 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way_status_out_81 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way_status_out_82 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way_status_out_83 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way_status_out_84 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way_status_out_85 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way_status_out_86 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way_status_out_87 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way_status_out_88 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way_status_out_89 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way_status_out_90 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way_status_out_91 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way_status_out_92 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way_status_out_93 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way_status_out_94 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way_status_out_95 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way_status_out_96 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way_status_out_97 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way_status_out_98 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way_status_out_99 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way_status_out_100 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way_status_out_101 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way_status_out_102 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way_status_out_103 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way_status_out_104 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way_status_out_105 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way_status_out_106 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way_status_out_107 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  way_status_out_108 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  way_status_out_109 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way_status_out_110 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way_status_out_111 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way_status_out_112 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way_status_out_113 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way_status_out_114 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way_status_out_115 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way_status_out_116 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way_status_out_117 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way_status_out_118 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way_status_out_119 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way_status_out_120 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way_status_out_121 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way_status_out_122 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way_status_out_123 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way_status_out_124 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way_status_out_125 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way_status_out_126 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way_status_out_127 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  tagv_mb_scnd_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_152[30:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  reset_ic_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  miss_addr = _RAND_160[25:0];
  _RAND_161 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_163[0:0];
  _RAND_164 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_164[63:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_441[0:0];
  _RAND_442 = {3{`RANDOM}};
  _T_1211 = _RAND_442[70:0];
  _RAND_443 = {1{`RANDOM}};
  ifc_region_acc_fault_memory_f = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_444[6:0];
  _RAND_445 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  bus_cmd_req_hold = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_448[2:0];
  _RAND_449 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_451[0:0];
  _RAND_452 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_452[38:0];
  _RAND_453 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_453[1:0];
  _RAND_454 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_454[2:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_dma_rtag_temp = _RAND_455[2:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_dma_rvalid_temp = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_dma_ecc_error = _RAND_457[0:0];
  _RAND_458 = {2{`RANDOM}};
  iccm_dma_rdata_temp = _RAND_458[63:0];
  _RAND_459 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_459[13:0];
  _RAND_460 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_461[13:0];
  _RAND_462 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_462[6:0];
  _RAND_463 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  way_status_new_ff = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_465[1:0];
  _RAND_466 = {1{`RANDOM}};
  ic_valid_ff = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_9798 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_9799 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_9800 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  _T_9804 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  _T_9805 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  _T_9826 = _RAND_472[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    flush_final_f = 1'h0;
  end
  if (reset) begin
    ifc_fetch_req_f_raw = 1'h0;
  end
  if (reset) begin
    miss_state = 3'h0;
  end
  if (reset) begin
    scnd_miss_req_q = 1'h0;
  end
  if (reset) begin
    ifu_fetch_addr_int_f = 31'h0;
  end
  if (reset) begin
    ifc_iccm_access_f = 1'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_in = 1'h0;
  end
  if (reset) begin
    dma_iccm_req_f = 1'h0;
  end
  if (reset) begin
    perr_state = 3'h0;
  end
  if (reset) begin
    err_stop_state = 2'h0;
  end
  if (reset) begin
    reset_all_tags = 1'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_final_f = 1'h0;
  end
  if (reset) begin
    ifu_bus_rvalid_unq_ff = 1'h0;
  end
  if (reset) begin
    bus_ifu_bus_clk_en_ff = 1'h0;
  end
  if (reset) begin
    uncacheable_miss_ff = 1'h0;
  end
  if (reset) begin
    bus_data_beat_count = 3'h0;
  end
  if (reset) begin
    ic_miss_buff_data_valid = 8'h0;
  end
  if (reset) begin
    imb_ff = 31'h0;
  end
  if (reset) begin
    last_data_recieved_ff = 1'h0;
  end
  if (reset) begin
    sel_mb_addr_ff = 1'h0;
  end
  if (reset) begin
    way_status_mb_scnd_ff = 1'h0;
  end
  if (reset) begin
    ifu_ic_rw_int_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_out_0 = 1'h0;
  end
  if (reset) begin
    way_status_out_1 = 1'h0;
  end
  if (reset) begin
    way_status_out_2 = 1'h0;
  end
  if (reset) begin
    way_status_out_3 = 1'h0;
  end
  if (reset) begin
    way_status_out_4 = 1'h0;
  end
  if (reset) begin
    way_status_out_5 = 1'h0;
  end
  if (reset) begin
    way_status_out_6 = 1'h0;
  end
  if (reset) begin
    way_status_out_7 = 1'h0;
  end
  if (reset) begin
    way_status_out_8 = 1'h0;
  end
  if (reset) begin
    way_status_out_9 = 1'h0;
  end
  if (reset) begin
    way_status_out_10 = 1'h0;
  end
  if (reset) begin
    way_status_out_11 = 1'h0;
  end
  if (reset) begin
    way_status_out_12 = 1'h0;
  end
  if (reset) begin
    way_status_out_13 = 1'h0;
  end
  if (reset) begin
    way_status_out_14 = 1'h0;
  end
  if (reset) begin
    way_status_out_15 = 1'h0;
  end
  if (reset) begin
    way_status_out_16 = 1'h0;
  end
  if (reset) begin
    way_status_out_17 = 1'h0;
  end
  if (reset) begin
    way_status_out_18 = 1'h0;
  end
  if (reset) begin
    way_status_out_19 = 1'h0;
  end
  if (reset) begin
    way_status_out_20 = 1'h0;
  end
  if (reset) begin
    way_status_out_21 = 1'h0;
  end
  if (reset) begin
    way_status_out_22 = 1'h0;
  end
  if (reset) begin
    way_status_out_23 = 1'h0;
  end
  if (reset) begin
    way_status_out_24 = 1'h0;
  end
  if (reset) begin
    way_status_out_25 = 1'h0;
  end
  if (reset) begin
    way_status_out_26 = 1'h0;
  end
  if (reset) begin
    way_status_out_27 = 1'h0;
  end
  if (reset) begin
    way_status_out_28 = 1'h0;
  end
  if (reset) begin
    way_status_out_29 = 1'h0;
  end
  if (reset) begin
    way_status_out_30 = 1'h0;
  end
  if (reset) begin
    way_status_out_31 = 1'h0;
  end
  if (reset) begin
    way_status_out_32 = 1'h0;
  end
  if (reset) begin
    way_status_out_33 = 1'h0;
  end
  if (reset) begin
    way_status_out_34 = 1'h0;
  end
  if (reset) begin
    way_status_out_35 = 1'h0;
  end
  if (reset) begin
    way_status_out_36 = 1'h0;
  end
  if (reset) begin
    way_status_out_37 = 1'h0;
  end
  if (reset) begin
    way_status_out_38 = 1'h0;
  end
  if (reset) begin
    way_status_out_39 = 1'h0;
  end
  if (reset) begin
    way_status_out_40 = 1'h0;
  end
  if (reset) begin
    way_status_out_41 = 1'h0;
  end
  if (reset) begin
    way_status_out_42 = 1'h0;
  end
  if (reset) begin
    way_status_out_43 = 1'h0;
  end
  if (reset) begin
    way_status_out_44 = 1'h0;
  end
  if (reset) begin
    way_status_out_45 = 1'h0;
  end
  if (reset) begin
    way_status_out_46 = 1'h0;
  end
  if (reset) begin
    way_status_out_47 = 1'h0;
  end
  if (reset) begin
    way_status_out_48 = 1'h0;
  end
  if (reset) begin
    way_status_out_49 = 1'h0;
  end
  if (reset) begin
    way_status_out_50 = 1'h0;
  end
  if (reset) begin
    way_status_out_51 = 1'h0;
  end
  if (reset) begin
    way_status_out_52 = 1'h0;
  end
  if (reset) begin
    way_status_out_53 = 1'h0;
  end
  if (reset) begin
    way_status_out_54 = 1'h0;
  end
  if (reset) begin
    way_status_out_55 = 1'h0;
  end
  if (reset) begin
    way_status_out_56 = 1'h0;
  end
  if (reset) begin
    way_status_out_57 = 1'h0;
  end
  if (reset) begin
    way_status_out_58 = 1'h0;
  end
  if (reset) begin
    way_status_out_59 = 1'h0;
  end
  if (reset) begin
    way_status_out_60 = 1'h0;
  end
  if (reset) begin
    way_status_out_61 = 1'h0;
  end
  if (reset) begin
    way_status_out_62 = 1'h0;
  end
  if (reset) begin
    way_status_out_63 = 1'h0;
  end
  if (reset) begin
    way_status_out_64 = 1'h0;
  end
  if (reset) begin
    way_status_out_65 = 1'h0;
  end
  if (reset) begin
    way_status_out_66 = 1'h0;
  end
  if (reset) begin
    way_status_out_67 = 1'h0;
  end
  if (reset) begin
    way_status_out_68 = 1'h0;
  end
  if (reset) begin
    way_status_out_69 = 1'h0;
  end
  if (reset) begin
    way_status_out_70 = 1'h0;
  end
  if (reset) begin
    way_status_out_71 = 1'h0;
  end
  if (reset) begin
    way_status_out_72 = 1'h0;
  end
  if (reset) begin
    way_status_out_73 = 1'h0;
  end
  if (reset) begin
    way_status_out_74 = 1'h0;
  end
  if (reset) begin
    way_status_out_75 = 1'h0;
  end
  if (reset) begin
    way_status_out_76 = 1'h0;
  end
  if (reset) begin
    way_status_out_77 = 1'h0;
  end
  if (reset) begin
    way_status_out_78 = 1'h0;
  end
  if (reset) begin
    way_status_out_79 = 1'h0;
  end
  if (reset) begin
    way_status_out_80 = 1'h0;
  end
  if (reset) begin
    way_status_out_81 = 1'h0;
  end
  if (reset) begin
    way_status_out_82 = 1'h0;
  end
  if (reset) begin
    way_status_out_83 = 1'h0;
  end
  if (reset) begin
    way_status_out_84 = 1'h0;
  end
  if (reset) begin
    way_status_out_85 = 1'h0;
  end
  if (reset) begin
    way_status_out_86 = 1'h0;
  end
  if (reset) begin
    way_status_out_87 = 1'h0;
  end
  if (reset) begin
    way_status_out_88 = 1'h0;
  end
  if (reset) begin
    way_status_out_89 = 1'h0;
  end
  if (reset) begin
    way_status_out_90 = 1'h0;
  end
  if (reset) begin
    way_status_out_91 = 1'h0;
  end
  if (reset) begin
    way_status_out_92 = 1'h0;
  end
  if (reset) begin
    way_status_out_93 = 1'h0;
  end
  if (reset) begin
    way_status_out_94 = 1'h0;
  end
  if (reset) begin
    way_status_out_95 = 1'h0;
  end
  if (reset) begin
    way_status_out_96 = 1'h0;
  end
  if (reset) begin
    way_status_out_97 = 1'h0;
  end
  if (reset) begin
    way_status_out_98 = 1'h0;
  end
  if (reset) begin
    way_status_out_99 = 1'h0;
  end
  if (reset) begin
    way_status_out_100 = 1'h0;
  end
  if (reset) begin
    way_status_out_101 = 1'h0;
  end
  if (reset) begin
    way_status_out_102 = 1'h0;
  end
  if (reset) begin
    way_status_out_103 = 1'h0;
  end
  if (reset) begin
    way_status_out_104 = 1'h0;
  end
  if (reset) begin
    way_status_out_105 = 1'h0;
  end
  if (reset) begin
    way_status_out_106 = 1'h0;
  end
  if (reset) begin
    way_status_out_107 = 1'h0;
  end
  if (reset) begin
    way_status_out_108 = 1'h0;
  end
  if (reset) begin
    way_status_out_109 = 1'h0;
  end
  if (reset) begin
    way_status_out_110 = 1'h0;
  end
  if (reset) begin
    way_status_out_111 = 1'h0;
  end
  if (reset) begin
    way_status_out_112 = 1'h0;
  end
  if (reset) begin
    way_status_out_113 = 1'h0;
  end
  if (reset) begin
    way_status_out_114 = 1'h0;
  end
  if (reset) begin
    way_status_out_115 = 1'h0;
  end
  if (reset) begin
    way_status_out_116 = 1'h0;
  end
  if (reset) begin
    way_status_out_117 = 1'h0;
  end
  if (reset) begin
    way_status_out_118 = 1'h0;
  end
  if (reset) begin
    way_status_out_119 = 1'h0;
  end
  if (reset) begin
    way_status_out_120 = 1'h0;
  end
  if (reset) begin
    way_status_out_121 = 1'h0;
  end
  if (reset) begin
    way_status_out_122 = 1'h0;
  end
  if (reset) begin
    way_status_out_123 = 1'h0;
  end
  if (reset) begin
    way_status_out_124 = 1'h0;
  end
  if (reset) begin
    way_status_out_125 = 1'h0;
  end
  if (reset) begin
    way_status_out_126 = 1'h0;
  end
  if (reset) begin
    way_status_out_127 = 1'h0;
  end
  if (reset) begin
    tagv_mb_scnd_ff = 2'h0;
  end
  if (reset) begin
    uncacheable_miss_scnd_ff = 1'h0;
  end
  if (reset) begin
    imb_scnd_ff = 31'h0;
  end
  if (reset) begin
    ifu_bus_rid_ff = 3'h0;
  end
  if (reset) begin
    ifu_bus_rresp_ff = 2'h0;
  end
  if (reset) begin
    ifu_wr_data_comb_err_ff = 1'h0;
  end
  if (reset) begin
    way_status_mb_ff = 1'h0;
  end
  if (reset) begin
    tagv_mb_ff = 2'h0;
  end
  if (reset) begin
    reset_ic_ff = 1'h0;
  end
  if (reset) begin
    fetch_uncacheable_ff = 1'h0;
  end
  if (reset) begin
    miss_addr = 26'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_f = 1'h0;
  end
  if (reset) begin
    bus_rd_addr_count = 3'h0;
  end
  if (reset) begin
    ic_act_miss_f_delayed = 1'h0;
  end
  if (reset) begin
    ifu_bus_rdata_ff = 64'h0;
  end
  if (reset) begin
    ic_miss_buff_data_0 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_1 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_2 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_3 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_4 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_5 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_6 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_7 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_8 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_9 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_10 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_11 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_12 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_13 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_14 = 32'h0;
  end
  if (reset) begin
    ic_miss_buff_data_15 = 32'h0;
  end
  if (reset) begin
    ic_crit_wd_rdy_new_ff = 1'h0;
  end
  if (reset) begin
    ic_miss_buff_data_error = 8'h0;
  end
  if (reset) begin
    ic_debug_ict_array_sel_ff = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_1_127 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_0 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_1 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_2 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_3 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_4 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_5 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_6 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_7 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_8 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_9 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_10 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_11 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_12 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_13 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_14 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_15 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_16 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_17 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_18 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_19 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_20 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_21 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_22 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_23 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_24 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_25 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_26 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_27 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_28 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_29 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_30 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_31 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_32 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_33 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_34 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_35 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_36 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_37 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_38 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_39 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_40 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_41 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_42 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_43 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_44 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_45 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_46 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_47 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_48 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_49 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_50 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_51 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_52 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_53 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_54 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_55 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_56 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_57 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_58 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_59 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_60 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_61 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_62 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_63 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_64 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_65 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_66 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_67 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_68 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_69 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_70 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_71 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_72 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_73 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_74 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_75 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_76 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_77 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_78 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_79 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_80 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_81 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_82 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_83 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_84 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_85 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_86 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_87 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_88 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_89 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_90 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_91 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_92 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_93 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_94 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_95 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_96 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_97 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_98 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_99 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_100 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_101 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_102 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_103 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_104 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_105 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_106 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_107 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_108 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_109 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_110 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_111 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_112 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_113 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_114 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_115 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_116 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_117 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_118 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_119 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_120 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_121 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_122 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_123 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_124 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_125 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_126 = 1'h0;
  end
  if (reset) begin
    ic_tag_valid_out_0_127 = 1'h0;
  end
  if (reset) begin
    ic_debug_way_ff = 2'h0;
  end
  if (reset) begin
    ic_debug_rd_en_ff = 1'h0;
  end
  if (reset) begin
    _T_1211 = 71'h0;
  end
  if (reset) begin
    ifc_region_acc_fault_memory_f = 1'h0;
  end
  if (reset) begin
    perr_ic_index_ff = 7'h0;
  end
  if (reset) begin
    dma_sb_err_state_ff = 1'h0;
  end
  if (reset) begin
    bus_cmd_req_hold = 1'h0;
  end
  if (reset) begin
    ifu_bus_cmd_valid = 1'h0;
  end
  if (reset) begin
    bus_cmd_beat_count = 3'h0;
  end
  if (reset) begin
    ifu_bus_arready_unq_ff = 1'h0;
  end
  if (reset) begin
    ifu_bus_arvalid_ff = 1'h0;
  end
  if (reset) begin
    ifc_dma_access_ok_prev = 1'h0;
  end
  if (reset) begin
    iccm_ecc_corr_data_ff = 39'h0;
  end
  if (reset) begin
    dma_mem_addr_ff = 2'h0;
  end
  if (reset) begin
    dma_mem_tag_ff = 3'h0;
  end
  if (reset) begin
    iccm_dma_rtag_temp = 3'h0;
  end
  if (reset) begin
    iccm_dma_rvalid_temp = 1'h0;
  end
  if (reset) begin
    iccm_dma_ecc_error = 1'h0;
  end
  if (reset) begin
    iccm_dma_rdata_temp = 64'h0;
  end
  if (reset) begin
    iccm_ecc_corr_index_ff = 14'h0;
  end
  if (reset) begin
    iccm_rd_ecc_single_err_ff = 1'h0;
  end
  if (reset) begin
    iccm_rw_addr_f = 14'h0;
  end
  if (reset) begin
    ifu_status_wr_addr_ff = 7'h0;
  end
  if (reset) begin
    way_status_wr_en_ff = 1'h0;
  end
  if (reset) begin
    way_status_new_ff = 1'h0;
  end
  if (reset) begin
    ifu_tag_wren_ff = 2'h0;
  end
  if (reset) begin
    ic_valid_ff = 1'h0;
  end
  if (reset) begin
    _T_9798 = 1'h0;
  end
  if (reset) begin
    _T_9799 = 1'h0;
  end
  if (reset) begin
    _T_9800 = 1'h0;
  end
  if (reset) begin
    _T_9804 = 1'h0;
  end
  if (reset) begin
    _T_9805 = 1'h0;
  end
  if (reset) begin
    _T_9826 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= _T_317 & _T_318;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= _T_22 & _T_319;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2708 & _T_2712;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2499) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2501) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2511) begin
        perr_state <= 3'h0;
      end else if (_T_2514) begin
        if (_T_2517) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2521) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2525) begin
        err_stop_state <= 2'h1;
      end else if (_T_2530) begin
        if (_T_2532) begin
          err_stop_state <= 2'h0;
        end else if (_T_2553) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2557) begin
        if (_T_2532) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2574) begin
        if (_T_2578) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf | ifc_region_acc_fault_memory_bf;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= _T_2630 | _T_2631;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= {_T_1357,ic_miss_buff_data_valid_in_0};
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      imb_ff <= 31'h0;
    end else if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= _T_2638 | _T_2640;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= _T_334 | reset_tag_valid_for_miss;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_ic_rw_int_addr_ff <= 7'h0;
    end else if (_T_3996) begin
      ifu_ic_rw_int_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_ic_rw_int_addr_ff <= ifu_ic_rw_int_addr[11:5];
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_0 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_0 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_1 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_1 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_2 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_2 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_3 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_3 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_4 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_4 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_5 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_5 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_6 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_6 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_70_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_7 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_7 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_8 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_8 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_9 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_9 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_10 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_10 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_11 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_11 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_12 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_12 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_13 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_13 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_14 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_14 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_71_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_15 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_15 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_16 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_16 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_17 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_17 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_18 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_18 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_19 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_19 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_20 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_20 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_21 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_21 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_22 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_22 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_72_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_23 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_23 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_24 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_24 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_25 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_25 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_26 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_26 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_27 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_27 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_28 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_28 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_29 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_29 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_30 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_30 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_73_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_31 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_31 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_32 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_32 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_33 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_33 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_34 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_34 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_35 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_35 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_36 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_36 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_37 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_37 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_38 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_38 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_74_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_39 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_39 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_40 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_40 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_41 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_41 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_42 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_42 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_43 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_43 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_44 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_44 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_45 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_45 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_46 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_46 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_75_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_47 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_47 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_48 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_48 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_49 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_49 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_50 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_50 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_51 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_51 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_52 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_52 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_53 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_53 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_54 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_54 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_76_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_55 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_55 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_56 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_56 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_57 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_57 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_58 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_58 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_59 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_59 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_60 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_60 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_61 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_61 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_62 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_62 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_77_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_63 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_63 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_64 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_64 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_65 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_65 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_66 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_66 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_67 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_67 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_68 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_68 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_69 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_69 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_70 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_70 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_78_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_71 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_71 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_72 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_72 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_73 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_73 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_74 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_74 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_75 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_75 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_76 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_76 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_77 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_77 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_78 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_78 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_79_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_79 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_79 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_80 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_80 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_81 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_81 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_82 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_82 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_83 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_83 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_84 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_84 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_85 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_85 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_86 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_86 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_80_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_87 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_87 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_88 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_88 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_89 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_89 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_90 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_90 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_91 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_91 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_92 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_92 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_93 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_93 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_94 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_94 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_81_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_95 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_95 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_96 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_96 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_97 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_97 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_98 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_98 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_99 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_99 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_100 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_100 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_101 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_101 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_102 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_102 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_82_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_103 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_103 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_104 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_104 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_105 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_105 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_106 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_106 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_107 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_107 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_108 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_108 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_109 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_109 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_110 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_110 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_83_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_111 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_111 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_112 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_112 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_113 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_113 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_114 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_114 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_115 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_115 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_116 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_116 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_117 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_117 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_118 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_118 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_84_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_119 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_119 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_120 <= 1'h0;
    end else if (_T_4020) begin
      way_status_out_120 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_121 <= 1'h0;
    end else if (_T_4024) begin
      way_status_out_121 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_122 <= 1'h0;
    end else if (_T_4028) begin
      way_status_out_122 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_123 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_123 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_124 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_124 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_125 <= 1'h0;
    end else if (_T_4040) begin
      way_status_out_125 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_126 <= 1'h0;
    end else if (_T_4044) begin
      way_status_out_126 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_85_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_out_127 <= 1'h0;
    end else if (_T_4048) begin
      way_status_out_127 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      tagv_mb_scnd_ff <= 2'h0;
    end else if (!(_T_19)) begin
      tagv_mb_scnd_ff <= _T_198;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err_data & _T_2626;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_290;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= _T_295;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      reset_ic_ff <= 1'h0;
    end else begin
      reset_ic_ff <= _T_298 & _T_299;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_231) begin
      bus_rd_addr_count <= imb_ff[4:2];
    end else if (scnd_miss_req_q) begin
      bus_rd_addr_count <= imb_scnd_ff[4:2];
    end else if (bus_cmd_sent) begin
      bus_rd_addr_count <= _T_2646;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= _T_233 & _T_209;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_31_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_40_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_40_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_49_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_49_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_58_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_58_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge rvclkhdr_67_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
  end
  always @(posedge rvclkhdr_67_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= _T_1513 | _T_1518;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= {_T_1397,ic_miss_buff_data_error_in_0};
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else begin
      ic_debug_ict_array_sel_ff <= io_ic_debug_rd_en & io_ic_debug_tag_array;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5641) begin
      ic_tag_valid_out_1_0 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5656) begin
      ic_tag_valid_out_1_1 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5671) begin
      ic_tag_valid_out_1_2 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5686) begin
      ic_tag_valid_out_1_3 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5701) begin
      ic_tag_valid_out_1_4 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5716) begin
      ic_tag_valid_out_1_5 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5731) begin
      ic_tag_valid_out_1_6 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5746) begin
      ic_tag_valid_out_1_7 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5761) begin
      ic_tag_valid_out_1_8 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5776) begin
      ic_tag_valid_out_1_9 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5791) begin
      ic_tag_valid_out_1_10 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5806) begin
      ic_tag_valid_out_1_11 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5821) begin
      ic_tag_valid_out_1_12 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5836) begin
      ic_tag_valid_out_1_13 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5851) begin
      ic_tag_valid_out_1_14 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5866) begin
      ic_tag_valid_out_1_15 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5881) begin
      ic_tag_valid_out_1_16 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5896) begin
      ic_tag_valid_out_1_17 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5911) begin
      ic_tag_valid_out_1_18 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5926) begin
      ic_tag_valid_out_1_19 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5941) begin
      ic_tag_valid_out_1_20 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5956) begin
      ic_tag_valid_out_1_21 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5971) begin
      ic_tag_valid_out_1_22 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5986) begin
      ic_tag_valid_out_1_23 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6001) begin
      ic_tag_valid_out_1_24 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6016) begin
      ic_tag_valid_out_1_25 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6031) begin
      ic_tag_valid_out_1_26 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6046) begin
      ic_tag_valid_out_1_27 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6061) begin
      ic_tag_valid_out_1_28 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6076) begin
      ic_tag_valid_out_1_29 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6091) begin
      ic_tag_valid_out_1_30 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_87_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6106) begin
      ic_tag_valid_out_1_31 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6601) begin
      ic_tag_valid_out_1_32 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6616) begin
      ic_tag_valid_out_1_33 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6631) begin
      ic_tag_valid_out_1_34 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6646) begin
      ic_tag_valid_out_1_35 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6661) begin
      ic_tag_valid_out_1_36 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6676) begin
      ic_tag_valid_out_1_37 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6691) begin
      ic_tag_valid_out_1_38 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6706) begin
      ic_tag_valid_out_1_39 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6721) begin
      ic_tag_valid_out_1_40 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6736) begin
      ic_tag_valid_out_1_41 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6751) begin
      ic_tag_valid_out_1_42 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6766) begin
      ic_tag_valid_out_1_43 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6781) begin
      ic_tag_valid_out_1_44 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6796) begin
      ic_tag_valid_out_1_45 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6811) begin
      ic_tag_valid_out_1_46 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6826) begin
      ic_tag_valid_out_1_47 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6841) begin
      ic_tag_valid_out_1_48 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6856) begin
      ic_tag_valid_out_1_49 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6871) begin
      ic_tag_valid_out_1_50 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6886) begin
      ic_tag_valid_out_1_51 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6901) begin
      ic_tag_valid_out_1_52 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6916) begin
      ic_tag_valid_out_1_53 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6931) begin
      ic_tag_valid_out_1_54 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6946) begin
      ic_tag_valid_out_1_55 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6961) begin
      ic_tag_valid_out_1_56 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6976) begin
      ic_tag_valid_out_1_57 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6991) begin
      ic_tag_valid_out_1_58 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7006) begin
      ic_tag_valid_out_1_59 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7021) begin
      ic_tag_valid_out_1_60 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7036) begin
      ic_tag_valid_out_1_61 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7051) begin
      ic_tag_valid_out_1_62 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_89_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7066) begin
      ic_tag_valid_out_1_63 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7561) begin
      ic_tag_valid_out_1_64 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7576) begin
      ic_tag_valid_out_1_65 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7591) begin
      ic_tag_valid_out_1_66 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7606) begin
      ic_tag_valid_out_1_67 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7621) begin
      ic_tag_valid_out_1_68 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7636) begin
      ic_tag_valid_out_1_69 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7651) begin
      ic_tag_valid_out_1_70 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7666) begin
      ic_tag_valid_out_1_71 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7681) begin
      ic_tag_valid_out_1_72 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7696) begin
      ic_tag_valid_out_1_73 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7711) begin
      ic_tag_valid_out_1_74 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7726) begin
      ic_tag_valid_out_1_75 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7741) begin
      ic_tag_valid_out_1_76 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7756) begin
      ic_tag_valid_out_1_77 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7771) begin
      ic_tag_valid_out_1_78 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7786) begin
      ic_tag_valid_out_1_79 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7801) begin
      ic_tag_valid_out_1_80 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7816) begin
      ic_tag_valid_out_1_81 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7831) begin
      ic_tag_valid_out_1_82 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7846) begin
      ic_tag_valid_out_1_83 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7861) begin
      ic_tag_valid_out_1_84 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7876) begin
      ic_tag_valid_out_1_85 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7891) begin
      ic_tag_valid_out_1_86 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7906) begin
      ic_tag_valid_out_1_87 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_7921) begin
      ic_tag_valid_out_1_88 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_7936) begin
      ic_tag_valid_out_1_89 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_7951) begin
      ic_tag_valid_out_1_90 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_7966) begin
      ic_tag_valid_out_1_91 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_7981) begin
      ic_tag_valid_out_1_92 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_7996) begin
      ic_tag_valid_out_1_93 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8011) begin
      ic_tag_valid_out_1_94 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_91_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8026) begin
      ic_tag_valid_out_1_95 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8521) begin
      ic_tag_valid_out_1_96 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8536) begin
      ic_tag_valid_out_1_97 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8551) begin
      ic_tag_valid_out_1_98 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8566) begin
      ic_tag_valid_out_1_99 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8581) begin
      ic_tag_valid_out_1_100 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8596) begin
      ic_tag_valid_out_1_101 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8611) begin
      ic_tag_valid_out_1_102 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8626) begin
      ic_tag_valid_out_1_103 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8641) begin
      ic_tag_valid_out_1_104 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8656) begin
      ic_tag_valid_out_1_105 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8671) begin
      ic_tag_valid_out_1_106 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8686) begin
      ic_tag_valid_out_1_107 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8701) begin
      ic_tag_valid_out_1_108 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8716) begin
      ic_tag_valid_out_1_109 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8731) begin
      ic_tag_valid_out_1_110 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8746) begin
      ic_tag_valid_out_1_111 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8761) begin
      ic_tag_valid_out_1_112 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8776) begin
      ic_tag_valid_out_1_113 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8791) begin
      ic_tag_valid_out_1_114 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_8806) begin
      ic_tag_valid_out_1_115 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_8821) begin
      ic_tag_valid_out_1_116 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_8836) begin
      ic_tag_valid_out_1_117 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_8851) begin
      ic_tag_valid_out_1_118 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_8866) begin
      ic_tag_valid_out_1_119 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_8881) begin
      ic_tag_valid_out_1_120 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_8896) begin
      ic_tag_valid_out_1_121 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_8911) begin
      ic_tag_valid_out_1_122 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_8926) begin
      ic_tag_valid_out_1_123 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_8941) begin
      ic_tag_valid_out_1_124 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_8956) begin
      ic_tag_valid_out_1_125 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_8971) begin
      ic_tag_valid_out_1_126 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_93_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_8986) begin
      ic_tag_valid_out_1_127 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5161) begin
      ic_tag_valid_out_0_0 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5176) begin
      ic_tag_valid_out_0_1 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5191) begin
      ic_tag_valid_out_0_2 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5206) begin
      ic_tag_valid_out_0_3 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5221) begin
      ic_tag_valid_out_0_4 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5236) begin
      ic_tag_valid_out_0_5 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5251) begin
      ic_tag_valid_out_0_6 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5266) begin
      ic_tag_valid_out_0_7 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5281) begin
      ic_tag_valid_out_0_8 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5296) begin
      ic_tag_valid_out_0_9 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5311) begin
      ic_tag_valid_out_0_10 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5326) begin
      ic_tag_valid_out_0_11 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5341) begin
      ic_tag_valid_out_0_12 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5356) begin
      ic_tag_valid_out_0_13 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5371) begin
      ic_tag_valid_out_0_14 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5386) begin
      ic_tag_valid_out_0_15 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5401) begin
      ic_tag_valid_out_0_16 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5416) begin
      ic_tag_valid_out_0_17 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5431) begin
      ic_tag_valid_out_0_18 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5446) begin
      ic_tag_valid_out_0_19 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5461) begin
      ic_tag_valid_out_0_20 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5476) begin
      ic_tag_valid_out_0_21 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5491) begin
      ic_tag_valid_out_0_22 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5506) begin
      ic_tag_valid_out_0_23 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5521) begin
      ic_tag_valid_out_0_24 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5536) begin
      ic_tag_valid_out_0_25 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5551) begin
      ic_tag_valid_out_0_26 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5566) begin
      ic_tag_valid_out_0_27 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5581) begin
      ic_tag_valid_out_0_28 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5596) begin
      ic_tag_valid_out_0_29 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5611) begin
      ic_tag_valid_out_0_30 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_86_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5626) begin
      ic_tag_valid_out_0_31 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6121) begin
      ic_tag_valid_out_0_32 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6136) begin
      ic_tag_valid_out_0_33 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6151) begin
      ic_tag_valid_out_0_34 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6166) begin
      ic_tag_valid_out_0_35 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6181) begin
      ic_tag_valid_out_0_36 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6196) begin
      ic_tag_valid_out_0_37 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6211) begin
      ic_tag_valid_out_0_38 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6226) begin
      ic_tag_valid_out_0_39 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6241) begin
      ic_tag_valid_out_0_40 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6256) begin
      ic_tag_valid_out_0_41 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6271) begin
      ic_tag_valid_out_0_42 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6286) begin
      ic_tag_valid_out_0_43 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6301) begin
      ic_tag_valid_out_0_44 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6316) begin
      ic_tag_valid_out_0_45 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6331) begin
      ic_tag_valid_out_0_46 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6346) begin
      ic_tag_valid_out_0_47 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6361) begin
      ic_tag_valid_out_0_48 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6376) begin
      ic_tag_valid_out_0_49 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6391) begin
      ic_tag_valid_out_0_50 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6406) begin
      ic_tag_valid_out_0_51 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6421) begin
      ic_tag_valid_out_0_52 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6436) begin
      ic_tag_valid_out_0_53 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6451) begin
      ic_tag_valid_out_0_54 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6466) begin
      ic_tag_valid_out_0_55 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6481) begin
      ic_tag_valid_out_0_56 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6496) begin
      ic_tag_valid_out_0_57 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6511) begin
      ic_tag_valid_out_0_58 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6526) begin
      ic_tag_valid_out_0_59 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6541) begin
      ic_tag_valid_out_0_60 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6556) begin
      ic_tag_valid_out_0_61 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6571) begin
      ic_tag_valid_out_0_62 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_88_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6586) begin
      ic_tag_valid_out_0_63 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7081) begin
      ic_tag_valid_out_0_64 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7096) begin
      ic_tag_valid_out_0_65 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7111) begin
      ic_tag_valid_out_0_66 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7126) begin
      ic_tag_valid_out_0_67 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7141) begin
      ic_tag_valid_out_0_68 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7156) begin
      ic_tag_valid_out_0_69 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7171) begin
      ic_tag_valid_out_0_70 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7186) begin
      ic_tag_valid_out_0_71 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7201) begin
      ic_tag_valid_out_0_72 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7216) begin
      ic_tag_valid_out_0_73 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7231) begin
      ic_tag_valid_out_0_74 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7246) begin
      ic_tag_valid_out_0_75 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7261) begin
      ic_tag_valid_out_0_76 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7276) begin
      ic_tag_valid_out_0_77 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7291) begin
      ic_tag_valid_out_0_78 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7306) begin
      ic_tag_valid_out_0_79 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7321) begin
      ic_tag_valid_out_0_80 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7336) begin
      ic_tag_valid_out_0_81 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7351) begin
      ic_tag_valid_out_0_82 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7366) begin
      ic_tag_valid_out_0_83 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7381) begin
      ic_tag_valid_out_0_84 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7396) begin
      ic_tag_valid_out_0_85 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7411) begin
      ic_tag_valid_out_0_86 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7426) begin
      ic_tag_valid_out_0_87 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7441) begin
      ic_tag_valid_out_0_88 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7456) begin
      ic_tag_valid_out_0_89 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7471) begin
      ic_tag_valid_out_0_90 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7486) begin
      ic_tag_valid_out_0_91 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7501) begin
      ic_tag_valid_out_0_92 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7516) begin
      ic_tag_valid_out_0_93 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7531) begin
      ic_tag_valid_out_0_94 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_90_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7546) begin
      ic_tag_valid_out_0_95 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8041) begin
      ic_tag_valid_out_0_96 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8056) begin
      ic_tag_valid_out_0_97 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8071) begin
      ic_tag_valid_out_0_98 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8086) begin
      ic_tag_valid_out_0_99 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8101) begin
      ic_tag_valid_out_0_100 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8116) begin
      ic_tag_valid_out_0_101 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8131) begin
      ic_tag_valid_out_0_102 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8146) begin
      ic_tag_valid_out_0_103 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8161) begin
      ic_tag_valid_out_0_104 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8176) begin
      ic_tag_valid_out_0_105 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8191) begin
      ic_tag_valid_out_0_106 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8206) begin
      ic_tag_valid_out_0_107 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8221) begin
      ic_tag_valid_out_0_108 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8236) begin
      ic_tag_valid_out_0_109 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8251) begin
      ic_tag_valid_out_0_110 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8266) begin
      ic_tag_valid_out_0_111 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8281) begin
      ic_tag_valid_out_0_112 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8296) begin
      ic_tag_valid_out_0_113 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8311) begin
      ic_tag_valid_out_0_114 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8326) begin
      ic_tag_valid_out_0_115 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8341) begin
      ic_tag_valid_out_0_116 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8356) begin
      ic_tag_valid_out_0_117 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8371) begin
      ic_tag_valid_out_0_118 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8386) begin
      ic_tag_valid_out_0_119 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8401) begin
      ic_tag_valid_out_0_120 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8416) begin
      ic_tag_valid_out_0_121 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8431) begin
      ic_tag_valid_out_0_122 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8446) begin
      ic_tag_valid_out_0_123 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8461) begin
      ic_tag_valid_out_0_124 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8476) begin
      ic_tag_valid_out_0_125 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8491) begin
      ic_tag_valid_out_0_126 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_92_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8506) begin
      ic_tag_valid_out_0_127 <= _T_5153;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk or posedge reset) begin
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
  end
  always @(posedge rvclkhdr_io_l1clk or posedge reset) begin
    if (reset) begin
      _T_1211 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1211 <= _T_1210;
    end else begin
      _T_1211 <= io_ic_debug_rd_data;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifc_region_acc_fault_memory_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_memory_f <= _T_9885 & io_ifc_fetch_req_bf;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      perr_ic_index_ff <= 7'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= perr_state == 3'h4;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      bus_cmd_req_hold <= 1'h0;
    end else begin
      bus_cmd_req_hold <= _T_2603 & _T_2622;
    end
  end
  always @(posedge rvclkhdr_69_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else begin
      ifu_bus_cmd_valid <= _T_2593 & _T_2599;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk or posedge reset) begin
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (bus_cmd_beat_en) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
  end
  always @(posedge rvclkhdr_68_io_l1clk or posedge reset) begin
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= _T_2698 & _T_2699;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3931;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rtag_temp <= 3'h0;
    end else begin
      iccm_dma_rtag_temp <= dma_mem_tag_ff;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rvalid_temp <= 1'h0;
    end else begin
      iccm_dma_rvalid_temp <= iccm_dma_rvalid_in;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_ecc_error <= 1'h0;
    end else begin
      iccm_dma_ecc_error <= |iccm_double_ecc_error;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_dma_rdata_temp <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata_temp <= _T_3103;
    end else begin
      iccm_dma_rdata_temp <= _T_3104;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3927;
      end
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= _T_3922 & _T_319;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3996) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en | _T_3999;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      way_status_new_ff <= 1'h0;
    end else if (_T_3999) begin
      way_status_new_ff <= io_ic_debug_wr_data[4];
    end else if (_T_9776) begin
      way_status_new_ff <= replace_way_mb_any_0;
    end else begin
      way_status_new_ff <= way_status_hit_new;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren | ic_debug_tag_wr_en;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3999) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9798 <= 1'h0;
    end else begin
      _T_9798 <= _T_233 & _T_209;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9799 <= 1'h0;
    end else begin
      _T_9799 <= _T_225 & _T_247;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9800 <= 1'h0;
    end else begin
      _T_9800 <= ic_byp_hit_f & ifu_byp_data_err_new;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9804 <= 1'h0;
    end else begin
      _T_9804 <= _T_9802 & miss_pending;
    end
  end
  always @(posedge io_active_clk or posedge reset) begin
    if (reset) begin
      _T_9805 <= 1'h0;
    end else begin
      _T_9805 <= _T_2617 & _T_2622;
    end
  end
  always @(posedge io_free_clk or posedge reset) begin
    if (reset) begin
      _T_9826 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_9826 <= ic_debug_rd_en_ff;
    end
  end
endmodule
